
module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         \u0/N46 , \u0/N45 , n1, n2, n3, n4, n5, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n579, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9434, n9435, n9436, n9437, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9474, n9475, n9476, n9477, n9569, n9570,
         n9571, n9572, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa23;
  wire   [7:0] sa13;
  wire   [7:0] sa03;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa22;
  wire   [7:0] sa12;
  wire   [7:0] sa02;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa21;
  wire   [7:0] sa11;
  wire   [7:0] sa01;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa20;
  wire   [7:0] sa10;
  wire   [7:0] sa00;
  wire   [31:0] \u0/rcon ;
  wire   [3:0] \u0/r0/rcnt ;
  assign text_in_r[127] = text_in[127];
  assign text_in_r[126] = text_in[126];
  assign text_in_r[125] = text_in[125];
  assign text_in_r[124] = text_in[124];
  assign text_in_r[123] = text_in[123];
  assign text_in_r[122] = text_in[122];
  assign text_in_r[121] = text_in[121];
  assign text_in_r[120] = text_in[120];
  assign text_in_r[119] = text_in[119];
  assign text_in_r[118] = text_in[118];
  assign text_in_r[117] = text_in[117];
  assign text_in_r[116] = text_in[116];
  assign text_in_r[115] = text_in[115];
  assign text_in_r[114] = text_in[114];
  assign text_in_r[113] = text_in[113];
  assign text_in_r[112] = text_in[112];
  assign text_in_r[111] = text_in[111];
  assign text_in_r[110] = text_in[110];
  assign text_in_r[109] = text_in[109];
  assign text_in_r[108] = text_in[108];
  assign text_in_r[107] = text_in[107];
  assign text_in_r[106] = text_in[106];
  assign text_in_r[105] = text_in[105];
  assign text_in_r[104] = text_in[104];
  assign text_in_r[103] = text_in[103];
  assign text_in_r[102] = text_in[102];
  assign text_in_r[101] = text_in[101];
  assign text_in_r[100] = text_in[100];
  assign text_in_r[99] = text_in[99];
  assign text_in_r[98] = text_in[98];
  assign text_in_r[97] = text_in[97];
  assign text_in_r[96] = text_in[96];
  assign text_in_r[95] = text_in[95];
  assign text_in_r[94] = text_in[94];
  assign text_in_r[93] = text_in[93];
  assign text_in_r[92] = text_in[92];
  assign text_in_r[91] = text_in[91];
  assign text_in_r[90] = text_in[90];
  assign text_in_r[89] = text_in[89];
  assign text_in_r[88] = text_in[88];
  assign text_in_r[87] = text_in[87];
  assign text_in_r[86] = text_in[86];
  assign text_in_r[85] = text_in[85];
  assign text_in_r[84] = text_in[84];
  assign text_in_r[83] = text_in[83];
  assign text_in_r[82] = text_in[82];
  assign text_in_r[81] = text_in[81];
  assign text_in_r[80] = text_in[80];
  assign text_in_r[79] = text_in[79];
  assign text_in_r[78] = text_in[78];
  assign text_in_r[77] = text_in[77];
  assign text_in_r[76] = text_in[76];
  assign text_in_r[75] = text_in[75];
  assign text_in_r[74] = text_in[74];
  assign text_in_r[73] = text_in[73];
  assign text_in_r[72] = text_in[72];
  assign text_in_r[71] = text_in[71];
  assign text_in_r[70] = text_in[70];
  assign text_in_r[69] = text_in[69];
  assign text_in_r[68] = text_in[68];
  assign text_in_r[67] = text_in[67];
  assign text_in_r[66] = text_in[66];
  assign text_in_r[65] = text_in[65];
  assign text_in_r[64] = text_in[64];
  assign text_in_r[63] = text_in[63];
  assign text_in_r[62] = text_in[62];
  assign text_in_r[61] = text_in[61];
  assign text_in_r[60] = text_in[60];
  assign text_in_r[59] = text_in[59];
  assign text_in_r[58] = text_in[58];
  assign text_in_r[57] = text_in[57];
  assign text_in_r[56] = text_in[56];
  assign text_in_r[55] = text_in[55];
  assign text_in_r[54] = text_in[54];
  assign text_in_r[53] = text_in[53];
  assign text_in_r[52] = text_in[52];
  assign text_in_r[51] = text_in[51];
  assign text_in_r[50] = text_in[50];
  assign text_in_r[49] = text_in[49];
  assign text_in_r[48] = text_in[48];
  assign text_in_r[47] = text_in[47];
  assign text_in_r[46] = text_in[46];
  assign text_in_r[45] = text_in[45];
  assign text_in_r[44] = text_in[44];
  assign text_in_r[43] = text_in[43];
  assign text_in_r[42] = text_in[42];
  assign text_in_r[41] = text_in[41];
  assign text_in_r[40] = text_in[40];
  assign text_in_r[39] = text_in[39];
  assign text_in_r[38] = text_in[38];
  assign text_in_r[37] = text_in[37];
  assign text_in_r[36] = text_in[36];
  assign text_in_r[35] = text_in[35];
  assign text_in_r[34] = text_in[34];
  assign text_in_r[33] = text_in[33];
  assign text_in_r[32] = text_in[32];
  assign text_in_r[31] = text_in[31];
  assign text_in_r[30] = text_in[30];
  assign text_in_r[29] = text_in[29];
  assign text_in_r[28] = text_in[28];
  assign text_in_r[27] = text_in[27];
  assign text_in_r[26] = text_in[26];
  assign text_in_r[25] = text_in[25];
  assign text_in_r[24] = text_in[24];
  assign text_in_r[23] = text_in[23];
  assign text_in_r[22] = text_in[22];
  assign text_in_r[21] = text_in[21];
  assign text_in_r[20] = text_in[20];
  assign text_in_r[19] = text_in[19];
  assign text_in_r[18] = text_in[18];
  assign text_in_r[17] = text_in[17];
  assign text_in_r[16] = text_in[16];
  assign text_in_r[15] = text_in[15];
  assign text_in_r[14] = text_in[14];
  assign text_in_r[13] = text_in[13];
  assign text_in_r[12] = text_in[12];
  assign text_in_r[11] = text_in[11];
  assign text_in_r[10] = text_in[10];
  assign text_in_r[9] = text_in[9];
  assign text_in_r[8] = text_in[8];
  assign text_in_r[7] = text_in[7];
  assign text_in_r[6] = text_in[6];
  assign text_in_r[5] = text_in[5];
  assign text_in_r[4] = text_in[4];
  assign text_in_r[3] = text_in[3];
  assign text_in_r[2] = text_in[2];
  assign text_in_r[1] = text_in[1];
  assign text_in_r[0] = text_in[0];

  HS65_LS_NOR4ABX2 U9553 ( .A(n4604), .B(n4605), .C(n4606), .D(n4607), .Z(
        n2831) );
  HS65_LS_NOR4ABX2 U9554 ( .A(n7980), .B(n7981), .C(n7982), .D(n7983), .Z(
        n2815) );
  HS65_LS_NOR4ABX2 U9555 ( .A(n6197), .B(n6198), .C(n6199), .D(n6200), .Z(
        n2823) );
  HS65_LS_NOR4ABX2 U9556 ( .A(n3900), .B(n3901), .C(n3902), .D(n3903), .Z(
        n2674) );
  HS65_LS_NOR4ABX2 U9557 ( .A(n8437), .B(n8438), .C(n8439), .D(n8440), .Z(
        n2813) );
  HS65_LS_NOR4ABX2 U9558 ( .A(n7876), .B(n7877), .C(n7878), .D(n7879), .Z(
        n2816) );
  HS65_LS_AND2X4 U9559 ( .A(n5751), .B(n5750), .Z(n4491) );
  HS65_LS_AND2X4 U9560 ( .A(n7343), .B(n7342), .Z(n6084) );
  HS65_LS_AND2X4 U9561 ( .A(n9058), .B(n9044), .Z(n7709) );
  HS65_LS_AND2X4 U9562 ( .A(n9116), .B(n9102), .Z(n7747) );
  HS65_LS_AND2X4 U9563 ( .A(n5813), .B(n5812), .Z(n4531) );
  HS65_LS_AND2X4 U9564 ( .A(n5946), .B(n5932), .Z(n4616) );
  HS65_LS_AND2X4 U9565 ( .A(n7538), .B(n7524), .Z(n6209) );
  HS65_LS_AND2X4 U9566 ( .A(n7479), .B(n7465), .Z(n6184) );
  HS65_LS_AND2X4 U9567 ( .A(n7405), .B(n7404), .Z(n6124) );
  HS65_LS_AND2X4 U9568 ( .A(n5887), .B(n5873), .Z(n4591) );
  HS65_LS_NOR2AX3 U9569 ( .A(n9385), .B(n469), .Z(n5924) );
  HS65_LS_NOR2AX3 U9570 ( .A(sa22[7]), .B(n250), .Z(n5865) );
  HS65_LS_NOR2AX3 U9571 ( .A(n9302), .B(n27), .Z(n5749) );
  HS65_LS_NOR2AX3 U9572 ( .A(n9390), .B(n292), .Z(n7516) );
  HS65_LS_NOR2AX3 U9573 ( .A(n9305), .B(n71), .Z(n7457) );
  HS65_LS_NOR2AX3 U9574 ( .A(n9381), .B(n553), .Z(n7341) );
  HS65_LS_NOR2AX3 U9575 ( .A(sa01[7]), .B(n509), .Z(n7403) );
  HS65_LS_NOR2AX3 U9576 ( .A(n9402), .B(n691), .Z(n5811) );
  HS65_LS_NOR2AX3 U9577 ( .A(sa20[1]), .B(n627), .Z(n9059) );
  HS65_LS_NOR2AX3 U9578 ( .A(n9241), .B(n140), .Z(n9117) );
  HS65_LS_NOR2AX3 U9579 ( .A(n9330), .B(n674), .Z(n4282) );
  HS65_LSS_XOR2X3 U9580 ( .A(n2727), .B(n2680), .Z(n2685) );
  HS65_LS_IVX2 U9581 ( .A(n4424), .Z(n451) );
  HS65_LS_IVX2 U9582 ( .A(n6017), .Z(n274) );
  HS65_LSS_XOR2X3 U9583 ( .A(n316), .B(n2761), .Z(n2629) );
  HS65_LSS_XOR2X3 U9584 ( .A(n2712), .B(n2660), .Z(n2666) );
  HS65_LSS_XNOR2X3 U9585 ( .A(n2828), .B(n2804), .Z(n4374) );
  HS65_LSS_XNOR2X3 U9586 ( .A(n2820), .B(n2796), .Z(n5967) );
  HS65_LSS_XNOR2X3 U9587 ( .A(n3223), .B(n2780), .Z(n4408) );
  HS65_LSS_XNOR2X3 U9588 ( .A(n3019), .B(n2772), .Z(n6001) );
  HS65_LSS_XOR2X3 U9589 ( .A(n2659), .B(n2668), .Z(n2711) );
  HS65_LSS_XOR2X3 U9590 ( .A(n2682), .B(n2687), .Z(n2725) );
  HS65_LSS_XOR2X3 U9591 ( .A(n3011), .B(n2764), .Z(n7592) );
  HS65_LS_IVX2 U9592 ( .A(n2908), .Z(n316) );
  HS65_LSS_XOR2X3 U9593 ( .A(n2812), .B(n7542), .Z(n7619) );
  HS65_LSS_XOR2X3 U9594 ( .A(n2828), .B(n4357), .Z(n4437) );
  HS65_LSS_XOR2X3 U9595 ( .A(n2820), .B(n5950), .Z(n6030) );
  HS65_LSS_XOR2X3 U9596 ( .A(n2712), .B(n2637), .Z(n2743) );
  HS65_LSS_XOR2X3 U9597 ( .A(n2660), .B(n2661), .Z(n2656) );
  HS65_LSS_XOR2X3 U9598 ( .A(n3011), .B(n7556), .Z(n7553) );
  HS65_LSS_XOR2X3 U9599 ( .A(n2727), .B(n2637), .Z(n2756) );
  HS65_LSS_XOR2X3 U9600 ( .A(n2680), .B(n2661), .Z(n2679) );
  HS65_LSS_XOR2X3 U9601 ( .A(n3019), .B(n274), .Z(n5961) );
  HS65_LSS_XOR2X3 U9602 ( .A(n3223), .B(n451), .Z(n4368) );
  HS65_LS_NOR3AX2 U9603 ( .A(n3029), .B(n3030), .C(n2919), .Z(n3025) );
  HS65_LS_NOR3AX2 U9604 ( .A(n2347), .B(n2358), .C(n2316), .Z(n2421) );
  HS65_LS_NOR3AX2 U9605 ( .A(n1595), .B(n1606), .C(n1564), .Z(n1669) );
  HS65_LS_NOR3AX2 U9606 ( .A(n1219), .B(n1230), .C(n1188), .Z(n1293) );
  HS65_LS_NOR3AX2 U9607 ( .A(n1971), .B(n1982), .C(n1940), .Z(n2045) );
  HS65_LS_NOR3AX2 U9608 ( .A(n8390), .B(n8401), .C(n8142), .Z(n8686) );
  HS65_LS_NOR3AX2 U9609 ( .A(n8450), .B(n8461), .C(n8174), .Z(n8774) );
  HS65_LS_NOR4ABX2 U9610 ( .A(n2251), .B(n2524), .C(n2516), .D(n2540), .Z(
        n2562) );
  HS65_LS_NOR4ABX2 U9611 ( .A(n1499), .B(n1772), .C(n1764), .D(n1788), .Z(
        n1810) );
  HS65_LS_NOR4ABX2 U9612 ( .A(n1875), .B(n2148), .C(n2140), .D(n2164), .Z(
        n2186) );
  HS65_LS_NOR4ABX2 U9613 ( .A(n1123), .B(n1396), .C(n1388), .D(n1412), .Z(
        n1434) );
  HS65_LS_NOR4ABX2 U9614 ( .A(n2888), .B(n3950), .C(n3960), .D(n4011), .Z(
        n4238) );
  HS65_LS_NOR4ABX2 U9615 ( .A(n3906), .B(n4060), .C(n4061), .D(n3934), .Z(
        n4056) );
  HS65_LS_NOR4ABX2 U9616 ( .A(n4090), .B(n4091), .C(n3924), .D(n3996), .Z(
        n4086) );
  HS65_LS_NOR4ABX2 U9617 ( .A(n2843), .B(n3971), .C(n3981), .D(n4035), .Z(
        n4297) );
  HS65_LS_NOR4ABX2 U9618 ( .A(n8347), .B(n7956), .C(n8337), .D(n8054), .Z(
        n8511) );
  HS65_LS_NOR4ABX2 U9619 ( .A(n4975), .B(n4953), .C(n4777), .D(n4612), .Z(
        n5367) );
  HS65_LS_NOR4ABX2 U9620 ( .A(n6568), .B(n6546), .C(n6370), .D(n6205), .Z(
        n6959) );
  HS65_LS_NOR4ABX2 U9621 ( .A(n6438), .B(n6415), .C(n6223), .D(n6135), .Z(
        n6726) );
  HS65_LS_NOR4ABX2 U9622 ( .A(n4845), .B(n4822), .C(n4630), .D(n4542), .Z(
        n5134) );
  HS65_LS_NOR4ABX2 U9623 ( .A(n95), .B(n8451), .C(n8175), .D(n7988), .Z(n8766)
         );
  HS65_LS_IVX2 U9624 ( .A(n8462), .Z(n95) );
  HS65_LS_NOR4ABX2 U9625 ( .A(n582), .B(n8391), .C(n8143), .D(n7975), .Z(n8678) );
  HS65_LS_IVX2 U9626 ( .A(n8402), .Z(n582) );
  HS65_LS_NOR4ABX2 U9627 ( .A(n2917), .B(n3029), .C(n3238), .D(n3248), .Z(
        n3550) );
  HS65_LS_NAND2X2 U9628 ( .A(n886), .B(n869), .Z(n1213) );
  HS65_LS_NAND2X2 U9629 ( .A(n927), .B(n910), .Z(n2341) );
  HS65_LS_NAND2X2 U9630 ( .A(n804), .B(n787), .Z(n1965) );
  HS65_LS_NAND2X2 U9631 ( .A(n845), .B(n828), .Z(n1589) );
  HS65_LS_NOR3AX2 U9632 ( .A(n3237), .B(n3249), .C(n3028), .Z(n3600) );
  HS65_LS_NOR3AX2 U9633 ( .A(n8336), .B(n8348), .C(n8053), .Z(n8545) );
  HS65_LS_NOR3AX2 U9634 ( .A(n3304), .B(n3316), .C(n3139), .Z(n3702) );
  HS65_LS_NOR3AX2 U9635 ( .A(n3075), .B(n3087), .C(n2936), .Z(n3459) );
  HS65_LS_NOR3AX2 U9636 ( .A(n8081), .B(n8105), .C(n8011), .Z(n8241) );
  HS65_LS_NOR4ABX2 U9637 ( .A(n6514), .B(n6492), .C(n6331), .D(n6193), .Z(
        n6842) );
  HS65_LS_NOR4ABX2 U9638 ( .A(n4921), .B(n4899), .C(n4738), .D(n4600), .Z(
        n5250) );
  HS65_LS_NOR4ABX2 U9639 ( .A(n6275), .B(n6298), .C(n6146), .D(n6079), .Z(
        n6603) );
  HS65_LS_NOR4ABX2 U9640 ( .A(n4682), .B(n4705), .C(n4553), .D(n4486), .Z(
        n5010) );
  HS65_LSS_XNOR2X3 U9641 ( .A(n2812), .B(n2788), .Z(n7560) );
  HS65_LS_IVX2 U9642 ( .A(n8411), .Z(n595) );
  HS65_LS_IVX2 U9643 ( .A(n8471), .Z(n108) );
  HS65_LS_IVX2 U9644 ( .A(n6646), .Z(n545) );
  HS65_LS_IVX2 U9645 ( .A(n5053), .Z(n19) );
  HS65_LS_IVX2 U9646 ( .A(n8562), .Z(n325) );
  HS65_LS_IVX4 U9653 ( .A(n9147), .Z(n9137) );
  HS65_LS_IVX4 U9654 ( .A(n9147), .Z(n9136) );
  HS65_LS_IVX2 U9655 ( .A(n9146), .Z(n9140) );
  HS65_LS_IVX2 U9656 ( .A(n9146), .Z(n9139) );
  HS65_LS_IVX2 U9657 ( .A(n9146), .Z(n9141) );
  HS65_LS_IVX2 U9658 ( .A(n9146), .Z(n9138) );
  HS65_LSS_XOR2X3 U9659 ( .A(n2768), .B(n2792), .Z(n7542) );
  HS65_LSS_XOR2X3 U9660 ( .A(n2808), .B(n2784), .Z(n4357) );
  HS65_LSS_XOR2X3 U9661 ( .A(n2800), .B(n2776), .Z(n5950) );
  HS65_LSS_XOR2X3 U9662 ( .A(n2732), .B(n2728), .Z(n2637) );
  HS65_LSS_XOR2X3 U9663 ( .A(n2639), .B(n2691), .Z(n2661) );
  HS65_LSS_XNOR2X3 U9664 ( .A(n3015), .B(n2816), .Z(n7556) );
  HS65_LS_NOR4ABX2 U9665 ( .A(n7749), .B(n7750), .C(n7751), .D(n7752), .Z(
        n2761) );
  HS65_LS_MX41X4 U9666 ( .D0(n365), .S0(n399), .D1(n402), .S1(n369), .D2(n370), 
        .S2(n390), .D3(n376), .S3(n401), .Z(n7751) );
  HS65_LS_MX41X4 U9667 ( .D0(n398), .S0(n371), .D1(n380), .S1(n386), .D2(n378), 
        .S2(n396), .D3(n373), .S3(n7753), .Z(n7752) );
  HS65_LS_NOR4ABX2 U9668 ( .A(n7754), .B(n7755), .C(n7756), .D(n7757), .Z(
        n7750) );
  HS65_LS_NOR4ABX2 U9669 ( .A(n5010), .B(n5011), .C(n5012), .D(n5013), .Z(
        n2780) );
  HS65_LS_MX41X4 U9670 ( .D0(n25), .S0(n43), .D1(n31), .S1(n26), .D2(n29), 
        .S2(n23), .D3(n24), .S3(n4571), .Z(n5013) );
  HS65_LS_MX41X4 U9671 ( .D0(n14), .S0(n47), .D1(n45), .S1(n22), .D2(n48), 
        .S2(n20), .D3(n21), .S3(n33), .Z(n5012) );
  HS65_LS_AOI212X2 U9672 ( .A(n41), .B(n5014), .C(n18), .D(n4726), .E(n5015), 
        .Z(n5011) );
  HS65_LS_NOR4ABX2 U9673 ( .A(n6603), .B(n6604), .C(n6605), .D(n6606), .Z(
        n2772) );
  HS65_LS_MX41X4 U9674 ( .D0(n551), .S0(n569), .D1(n557), .S1(n552), .D2(n555), 
        .S2(n549), .D3(n550), .S3(n6164), .Z(n6606) );
  HS65_LS_MX41X4 U9675 ( .D0(n540), .S0(n573), .D1(n571), .S1(n548), .D2(n574), 
        .S2(n546), .D3(n547), .S3(n559), .Z(n6605) );
  HS65_LS_AOI212X2 U9676 ( .A(n567), .B(n6607), .C(n544), .D(n6319), .E(n6608), 
        .Z(n6604) );
  HS65_LS_NOR4ABX2 U9677 ( .A(n6842), .B(n6843), .C(n6844), .D(n6845), .Z(
        n2796) );
  HS65_LS_MX41X4 U9678 ( .D0(n63), .S0(n73), .D1(n77), .S1(n62), .D2(n74), 
        .S2(n59), .D3(n61), .S3(n80), .Z(n6844) );
  HS65_LS_MX41X4 U9679 ( .D0(n57), .S0(n87), .D1(n82), .S1(n58), .D2(n81), 
        .S2(n55), .D3(n56), .S3(n6348), .Z(n6845) );
  HS65_LS_AOI212X2 U9680 ( .A(n88), .B(n6846), .C(n60), .D(n6533), .E(n6847), 
        .Z(n6843) );
  HS65_LS_NOR4ABX2 U9681 ( .A(n5250), .B(n5251), .C(n5252), .D(n5253), .Z(
        n2804) );
  HS65_LS_MX41X4 U9682 ( .D0(n242), .S0(n252), .D1(n256), .S1(n241), .D2(n253), 
        .S2(n238), .D3(n240), .S3(n259), .Z(n5252) );
  HS65_LS_MX41X4 U9683 ( .D0(n236), .S0(n266), .D1(n261), .S1(n237), .D2(n260), 
        .S2(n234), .D3(n235), .S3(n4755), .Z(n5253) );
  HS65_LS_AOI212X2 U9684 ( .A(n267), .B(n5254), .C(n239), .D(n4940), .E(n5255), 
        .Z(n5251) );
  HS65_LS_NAND4ABX3 U9685 ( .A(n4295), .B(n4296), .C(n4297), .D(n4298), .Z(
        n2727) );
  HS65_LS_MX41X4 U9686 ( .D0(n440), .S0(n420), .D1(n431), .S1(n414), .D2(n415), 
        .S2(n441), .D3(n421), .S3(n3194), .Z(n4296) );
  HS65_LS_NOR4ABX2 U9687 ( .A(n3192), .B(n3844), .C(n4299), .D(n3858), .Z(
        n4298) );
  HS65_LS_MX41X4 U9688 ( .D0(n423), .S0(n439), .D1(n424), .S1(n435), .D2(n419), 
        .S2(n430), .D3(n410), .S3(n436), .Z(n4295) );
  HS65_LS_NAND4ABX3 U9689 ( .A(n4236), .B(n4237), .C(n4238), .D(n4239), .Z(
        n2680) );
  HS65_LS_MX41X4 U9690 ( .D0(n647), .S0(n663), .D1(n648), .S1(n659), .D2(n643), 
        .S2(n654), .D3(n633), .S3(n660), .Z(n4236) );
  HS65_LS_MX41X4 U9691 ( .D0(n664), .S0(n644), .D1(n655), .S1(n637), .D2(n639), 
        .S2(n665), .D3(n645), .S3(n3153), .Z(n4237) );
  HS65_LS_NOR4ABX2 U9692 ( .A(n3151), .B(n3727), .C(n4240), .D(n3741), .Z(
        n4239) );
  HS65_LS_NAND4ABX3 U9693 ( .A(n8764), .B(n8765), .C(n8766), .D(n8767), .Z(
        n2812) );
  HS65_LS_MX41X4 U9694 ( .D0(n98), .S0(n124), .D1(n119), .S1(n111), .D2(n113), 
        .S2(n122), .D3(n135), .S3(n114), .Z(n8764) );
  HS65_LS_MX41X4 U9695 ( .D0(n106), .S0(n133), .D1(n109), .S1(n137), .D2(n136), 
        .S2(n110), .D3(n107), .S3(n7748), .Z(n8765) );
  HS65_LS_AOI212X2 U9696 ( .A(n132), .B(n8768), .C(n112), .D(n7940), .E(n100), 
        .Z(n8767) );
  HS65_LS_NAND4ABX3 U9697 ( .A(n3783), .B(n3784), .C(n3785), .D(n3786), .Z(
        n2712) );
  HS65_LS_AOI212X2 U9698 ( .A(n446), .B(n3787), .C(n412), .D(n3395), .E(n3788), 
        .Z(n3786) );
  HS65_LS_MX41X4 U9699 ( .D0(n447), .S0(n417), .D1(n416), .S1(n437), .D2(n438), 
        .S2(n414), .D3(n415), .S3(n3194), .Z(n3784) );
  HS65_LS_MX41X4 U9700 ( .D0(n419), .S0(n430), .D1(n413), .S1(n434), .D2(n410), 
        .S2(n431), .D3(n436), .S3(n411), .Z(n3783) );
  HS65_LSS_XOR2X3 U9701 ( .A(n2832), .B(n2808), .Z(n4402) );
  HS65_LSS_XOR2X3 U9702 ( .A(n2824), .B(n2800), .Z(n5995) );
  HS65_LS_NAND4ABX3 U9703 ( .A(n6724), .B(n6725), .C(n6726), .D(n6727), .Z(
        n3019) );
  HS65_LS_MX41X4 U9704 ( .D0(n497), .S0(n529), .D1(n527), .S1(n504), .D2(n530), 
        .S2(n502), .D3(n503), .S3(n515), .Z(n6724) );
  HS65_LS_MX41X4 U9705 ( .D0(n507), .S0(n525), .D1(n513), .S1(n508), .D2(n511), 
        .S2(n505), .D3(n506), .S3(n6241), .Z(n6725) );
  HS65_LS_AOI212X2 U9706 ( .A(n523), .B(n6728), .C(n501), .D(n6459), .E(n6729), 
        .Z(n6727) );
  HS65_LS_NAND4ABX3 U9707 ( .A(n8509), .B(n8510), .C(n8511), .D(n8512), .Z(
        n3011) );
  HS65_LS_MX41X4 U9708 ( .D0(n335), .S0(n349), .D1(n326), .S1(n348), .D2(n323), 
        .S2(n346), .D3(n344), .S3(n327), .Z(n8509) );
  HS65_LS_MX41X4 U9709 ( .D0(n358), .S0(n332), .D1(n330), .S1(n345), .D2(n341), 
        .S2(n331), .D3(n329), .S3(n7784), .Z(n8510) );
  HS65_LS_AOI212X2 U9710 ( .A(n356), .B(n8513), .C(n324), .D(n8365), .E(n328), 
        .Z(n8512) );
  HS65_LS_NAND4ABX3 U9711 ( .A(n5365), .B(n5366), .C(n5367), .D(n5368), .Z(
        n2828) );
  HS65_LS_MX41X4 U9712 ( .D0(n461), .S0(n471), .D1(n475), .S1(n460), .D2(n472), 
        .S2(n457), .D3(n459), .S3(n478), .Z(n5365) );
  HS65_LS_MX41X4 U9713 ( .D0(n455), .S0(n485), .D1(n480), .S1(n456), .D2(n479), 
        .S2(n453), .D3(n454), .S3(n4794), .Z(n5366) );
  HS65_LS_AOI212X2 U9714 ( .A(n486), .B(n5369), .C(n458), .D(n4994), .E(n5370), 
        .Z(n5368) );
  HS65_LS_NAND4ABX3 U9715 ( .A(n6957), .B(n6958), .C(n6959), .D(n6960), .Z(
        n2820) );
  HS65_LS_MX41X4 U9716 ( .D0(n284), .S0(n294), .D1(n298), .S1(n283), .D2(n295), 
        .S2(n280), .D3(n282), .S3(n301), .Z(n6957) );
  HS65_LS_MX41X4 U9717 ( .D0(n278), .S0(n308), .D1(n303), .S1(n279), .D2(n302), 
        .S2(n276), .D3(n277), .S3(n6387), .Z(n6958) );
  HS65_LS_AOI212X2 U9718 ( .A(n309), .B(n6961), .C(n281), .D(n6587), .E(n6962), 
        .Z(n6960) );
  HS65_LS_NAND4ABX3 U9719 ( .A(n5132), .B(n5133), .C(n5134), .D(n5135), .Z(
        n3223) );
  HS65_LS_MX41X4 U9720 ( .D0(n679), .S0(n711), .D1(n709), .S1(n686), .D2(n712), 
        .S2(n684), .D3(n685), .S3(n697), .Z(n5132) );
  HS65_LS_MX41X4 U9721 ( .D0(n689), .S0(n707), .D1(n695), .S1(n690), .D2(n693), 
        .S2(n687), .D3(n688), .S3(n4648), .Z(n5133) );
  HS65_LS_AOI212X2 U9722 ( .A(n705), .B(n5136), .C(n683), .D(n4866), .E(n5137), 
        .Z(n5135) );
  HS65_LSS_XNOR2X3 U9723 ( .A(n2816), .B(n2792), .Z(n7586) );
  HS65_LSS_XOR2X3 U9724 ( .A(n3544), .B(n2784), .Z(n4813) );
  HS65_LSS_XOR2X3 U9725 ( .A(n3219), .B(n2776), .Z(n6406) );
  HS65_LS_NAND4ABX3 U9726 ( .A(n3666), .B(n3667), .C(n3668), .D(n3669), .Z(
        n2660) );
  HS65_LS_MX41X4 U9727 ( .D0(n671), .S0(n641), .D1(n640), .S1(n661), .D2(n662), 
        .S2(n637), .D3(n639), .S3(n3153), .Z(n3667) );
  HS65_LS_MX41X4 U9728 ( .D0(n643), .S0(n654), .D1(n636), .S1(n658), .D2(n633), 
        .S2(n655), .D3(n660), .S3(n634), .Z(n3666) );
  HS65_LS_AOI212X2 U9729 ( .A(n670), .B(n3670), .C(n635), .D(n3333), .E(n638), 
        .Z(n3669) );
  HS65_LSS_XOR2X3 U9730 ( .A(n2732), .B(n2691), .Z(n3229) );
  HS65_LS_NAND4ABX3 U9731 ( .A(n4084), .B(n4085), .C(n4086), .D(n4087), .Z(
        n2682) );
  HS65_LS_NOR4ABX2 U9732 ( .A(n3039), .B(n4088), .C(n3627), .D(n3642), .Z(
        n4087) );
  HS65_LS_MX41X4 U9733 ( .D0(n172), .S0(n152), .D1(n182), .S1(n153), .D2(n154), 
        .S2(n170), .D3(n150), .S3(n3050), .Z(n4085) );
  HS65_LS_MX41X4 U9734 ( .D0(n147), .S0(n171), .D1(n143), .S1(n167), .D2(n148), 
        .S2(n181), .D3(n158), .S3(n168), .Z(n4084) );
  HS65_LSS_XNOR2X3 U9735 ( .A(n2768), .B(n317), .Z(n2626) );
  HS65_LSS_XOR2X3 U9736 ( .A(n2815), .B(n2791), .Z(n7545) );
  HS65_LSS_XNOR2X3 U9737 ( .A(n2813), .B(n2789), .Z(n7554) );
  HS65_LS_NAND4ABX3 U9738 ( .A(n3548), .B(n3549), .C(n3550), .D(n3551), .Z(
        n2659) );
  HS65_LS_MX41X4 U9739 ( .D0(n177), .S0(n155), .D1(n156), .S1(n166), .D2(n165), 
        .S2(n153), .D3(n154), .S3(n3050), .Z(n3549) );
  HS65_LS_MX41X4 U9740 ( .D0(n148), .S0(n181), .D1(n159), .S1(n179), .D2(n158), 
        .S2(n182), .D3(n160), .S3(n168), .Z(n3548) );
  HS65_LS_AOI212X2 U9741 ( .A(n175), .B(n3552), .C(n157), .D(n3268), .E(n151), 
        .Z(n3551) );
  HS65_LS_NAND4ABX3 U9742 ( .A(n3422), .B(n3423), .C(n3424), .D(n3425), .Z(
        n2668) );
  HS65_LS_MX41X4 U9743 ( .D0(n193), .S0(n227), .D1(n204), .S1(n225), .D2(n203), 
        .S2(n228), .D3(n214), .S3(n205), .Z(n3422) );
  HS65_LS_MX41X4 U9744 ( .D0(n222), .S0(n200), .D1(n201), .S1(n212), .D2(n210), 
        .S2(n198), .D3(n199), .S3(n2951), .Z(n3423) );
  HS65_LS_AOI212X2 U9745 ( .A(n221), .B(n3426), .C(n202), .D(n3106), .E(n196), 
        .Z(n3425) );
  HS65_LSS_XOR2X3 U9746 ( .A(n2831), .B(n232), .Z(n4361) );
  HS65_LSS_XOR2X3 U9747 ( .A(n2823), .B(n52), .Z(n5954) );
  HS65_LSS_XOR2X3 U9748 ( .A(n2825), .B(n2801), .Z(n4387) );
  HS65_LSS_XOR2X3 U9749 ( .A(n2817), .B(n2793), .Z(n5980) );
  HS65_LSS_XOR2X3 U9750 ( .A(n3012), .B(n364), .Z(n7588) );
  HS65_LSS_XOR2X3 U9751 ( .A(n2707), .B(n2745), .Z(n2657) );
  HS65_LSS_XOR2X3 U9752 ( .A(n2809), .B(n2785), .Z(n2633) );
  HS65_LSS_XNOR2X3 U9753 ( .A(n3218), .B(n2775), .Z(n5987) );
  HS65_LSS_XNOR2X3 U9754 ( .A(n3220), .B(n2777), .Z(n4419) );
  HS65_LSS_XNOR2X3 U9755 ( .A(n3016), .B(n2769), .Z(n6012) );
  HS65_LSS_XNOR2X3 U9756 ( .A(n3543), .B(n2783), .Z(n4394) );
  HS65_LSS_XNOR2X3 U9757 ( .A(n3014), .B(n2767), .Z(n7578) );
  HS65_LS_NAND4ABX3 U9758 ( .A(n8204), .B(n8205), .C(n8206), .D(n8207), .Z(
        n2764) );
  HS65_LS_MX41X4 U9759 ( .D0(n395), .S0(n381), .D1(n379), .S1(n404), .D2(n403), 
        .S2(n380), .D3(n378), .S3(n7753), .Z(n8205) );
  HS65_LS_MX41X4 U9760 ( .D0(n370), .S0(n390), .D1(n377), .S1(n388), .D2(n376), 
        .S2(n386), .D3(n401), .S3(n375), .Z(n8204) );
  HS65_LS_AOI212X2 U9761 ( .A(n394), .B(n8208), .C(n374), .D(n8123), .E(n8209), 
        .Z(n8207) );
  HS65_LSS_XNOR2X3 U9762 ( .A(n2829), .B(n2805), .Z(n4369) );
  HS65_LSS_XOR2X3 U9763 ( .A(n2717), .B(n2667), .Z(n2673) );
  HS65_LS_NAND4ABX3 U9764 ( .A(n4054), .B(n4055), .C(n4056), .D(n4057), .Z(
        n2687) );
  HS65_LS_NOR4ABX2 U9765 ( .A(n2949), .B(n3485), .C(n4058), .D(n3500), .Z(
        n4057) );
  HS65_LS_MX41X4 U9766 ( .D0(n192), .S0(n218), .D1(n189), .S1(n213), .D2(n193), 
        .S2(n227), .D3(n203), .S3(n214), .Z(n4054) );
  HS65_LS_MX41X4 U9767 ( .D0(n217), .S0(n197), .D1(n228), .S1(n198), .D2(n199), 
        .S2(n216), .D3(n195), .S3(n2951), .Z(n4055) );
  HS65_LSS_XNOR2X3 U9768 ( .A(n2821), .B(n2797), .Z(n5962) );
  HS65_LSS_XOR2X3 U9769 ( .A(n2830), .B(n2806), .Z(n4365) );
  HS65_LSS_XOR2X3 U9770 ( .A(n2701), .B(n2647), .Z(n2651) );
  HS65_LSS_XNOR2X3 U9771 ( .A(n3224), .B(n2781), .Z(n4404) );
  HS65_LSS_XNOR2X3 U9772 ( .A(n2762), .B(n2630), .Z(n7600) );
  HS65_LSS_XNOR2X3 U9773 ( .A(n3216), .B(n2773), .Z(n5997) );
  HS65_LSS_XOR2X3 U9774 ( .A(n3010), .B(n362), .Z(n7595) );
  HS65_LSS_XNOR2X3 U9775 ( .A(n3013), .B(n2766), .Z(n7582) );
  HS65_LS_NAND4ABX3 U9776 ( .A(n8676), .B(n8677), .C(n8678), .D(n8679), .Z(
        n2788) );
  HS65_LS_MX41X4 U9777 ( .D0(n585), .S0(n611), .D1(n606), .S1(n598), .D2(n600), 
        .S2(n609), .D3(n622), .S3(n601), .Z(n8676) );
  HS65_LS_MX41X4 U9778 ( .D0(n593), .S0(n620), .D1(n596), .S1(n624), .D2(n623), 
        .S2(n597), .D3(n594), .S3(n7710), .Z(n8677) );
  HS65_LS_AOI212X2 U9779 ( .A(n619), .B(n8680), .C(n599), .D(n7841), .E(n587), 
        .Z(n8679) );
  HS65_LS_IVX2 U9780 ( .A(n2878), .Z(n199) );
  HS65_LSS_XNOR2X3 U9781 ( .A(n2674), .B(n2669), .Z(n2715) );
  HS65_LS_IVX2 U9782 ( .A(n7862), .Z(n378) );
  HS65_LSS_XNOR2X3 U9783 ( .A(n2818), .B(n51), .Z(n5975) );
  HS65_LSS_XNOR2X3 U9784 ( .A(n2722), .B(n629), .Z(n2677) );
  HS65_LSS_XNOR2X3 U9785 ( .A(n2646), .B(n186), .Z(n2699) );
  HS65_LSS_XNOR2X3 U9786 ( .A(n2640), .B(n188), .Z(n2694) );
  HS65_LSS_XNOR2X3 U9787 ( .A(n2653), .B(n187), .Z(n2706) );
  HS65_LSS_XNOR2X3 U9788 ( .A(n2681), .B(n142), .Z(n2721) );
  HS65_LS_AOI222X2 U9789 ( .A(n419), .B(n443), .C(n412), .D(n435), .E(n422), 
        .F(n446), .Z(n3810) );
  HS65_LSS_XNOR2X3 U9790 ( .A(n2827), .B(n233), .Z(n4379) );
  HS65_LSS_XNOR2X3 U9791 ( .A(n2819), .B(n53), .Z(n5972) );
  HS65_LSS_XNOR2X3 U9792 ( .A(n2696), .B(n631), .Z(n2644) );
  HS65_LSS_XNOR2X3 U9793 ( .A(n2811), .B(n577), .Z(n7565) );
  HS65_LS_NAND3X2 U9794 ( .A(n5715), .B(n5716), .C(n5717), .Z(n5514) );
  HS65_LS_NOR3AX2 U9795 ( .A(n4715), .B(n5081), .C(n5065), .Z(n5716) );
  HS65_LS_NOR3X1 U9796 ( .A(n5721), .B(n5043), .C(n5113), .Z(n5715) );
  HS65_LS_AOI212X2 U9797 ( .A(n17), .B(n33), .C(n15), .D(n46), .E(n5718), .Z(
        n5717) );
  HS65_LS_NAND3X2 U9798 ( .A(n7307), .B(n7308), .C(n7309), .Z(n7106) );
  HS65_LS_NOR3AX2 U9799 ( .A(n6308), .B(n6674), .C(n6658), .Z(n7308) );
  HS65_LS_NOR3X1 U9800 ( .A(n7313), .B(n6636), .C(n6706), .Z(n7307) );
  HS65_LS_AOI212X2 U9801 ( .A(n543), .B(n559), .C(n541), .D(n572), .E(n7310), 
        .Z(n7309) );
  HS65_LS_AOI222X2 U9802 ( .A(n210), .B(n189), .C(n217), .D(n199), .E(n212), 
        .F(n204), .Z(n4071) );
  HS65_LS_NAND4ABX3 U9803 ( .A(n1763), .B(n1764), .C(n1765), .D(n1766), .Z(
        n1761) );
  HS65_LS_AOI212X2 U9804 ( .A(n838), .B(n812), .C(n848), .D(n816), .E(n1500), 
        .Z(n1766) );
  HS65_LS_NAND4ABX3 U9805 ( .A(n2515), .B(n2516), .C(n2517), .D(n2518), .Z(
        n2513) );
  HS65_LS_AOI212X2 U9806 ( .A(n920), .B(n894), .C(n930), .D(n898), .E(n2252), 
        .Z(n2518) );
  HS65_LSS_XNOR2X3 U9807 ( .A(n2814), .B(n579), .Z(n7550) );
  HS65_LS_IVX2 U9808 ( .A(n2264), .Z(n910) );
  HS65_LS_IVX2 U9809 ( .A(n1136), .Z(n869) );
  HS65_LS_IVX2 U9810 ( .A(n1888), .Z(n787) );
  HS65_LS_IVX2 U9811 ( .A(n1512), .Z(n828) );
  HS65_LS_NAND3X2 U9812 ( .A(n8911), .B(n8912), .C(n8913), .Z(n8633) );
  HS65_LS_NOR3X1 U9813 ( .A(n8608), .B(n8359), .C(n8585), .Z(n8912) );
  HS65_LS_NOR3AX2 U9814 ( .A(n8623), .B(n8919), .C(n8568), .Z(n8911) );
  HS65_LS_AOI212X2 U9815 ( .A(n344), .B(n336), .C(n334), .D(n347), .E(n8914), 
        .Z(n8913) );
  HS65_LS_NAND3X2 U9816 ( .A(n4122), .B(n4123), .C(n4124), .Z(n3995) );
  HS65_LS_NOR3AX2 U9817 ( .A(n3565), .B(n4128), .C(n3256), .Z(n4122) );
  HS65_LS_NOR3AX2 U9818 ( .A(n3639), .B(n3655), .C(n3626), .Z(n4123) );
  HS65_LS_AOI212X2 U9819 ( .A(n168), .B(n150), .C(n149), .D(n180), .E(n4125), 
        .Z(n4124) );
  HS65_LS_AOI212X2 U9820 ( .A(n337), .B(n8553), .C(n330), .D(n354), .E(n8638), 
        .Z(n8637) );
  HS65_LS_CB4I6X4 U9821 ( .A(n324), .B(n329), .C(n348), .D(n8536), .Z(n8638)
         );
  HS65_LS_AOI212X2 U9822 ( .A(n371), .B(n8249), .C(n379), .D(n391), .E(n8670), 
        .Z(n8669) );
  HS65_LS_CB4I6X4 U9823 ( .A(n374), .B(n378), .C(n388), .D(n8319), .Z(n8670)
         );
  HS65_LS_AOI212X2 U9824 ( .A(n197), .B(n3467), .C(n201), .D(n223), .E(n4195), 
        .Z(n4194) );
  HS65_LS_CB4I6X4 U9825 ( .A(n202), .B(n199), .C(n225), .D(n3541), .Z(n4195)
         );
  HS65_LS_AOI212X2 U9826 ( .A(n928), .B(n894), .C(n925), .D(n906), .E(n2280), 
        .Z(n2273) );
  HS65_LS_OA12X4 U9827 ( .A(n2260), .B(n926), .C(n900), .Z(n2280) );
  HS65_LS_AOI212X2 U9828 ( .A(n846), .B(n812), .C(n843), .D(n824), .E(n1528), 
        .Z(n1521) );
  HS65_LS_OA12X4 U9829 ( .A(n1508), .B(n844), .C(n818), .Z(n1528) );
  HS65_LS_AOI222X2 U9830 ( .A(n780), .B(n794), .C(n776), .D(n806), .E(n792), 
        .F(n783), .Z(n2222) );
  HS65_LS_AOI222X2 U9831 ( .A(n862), .B(n876), .C(n858), .D(n888), .E(n874), 
        .F(n865), .Z(n1470) );
  HS65_LS_AOI222X2 U9832 ( .A(n399), .B(n367), .C(n401), .D(n375), .E(n376), 
        .F(n391), .Z(n8659) );
  HS65_LS_AOI222X2 U9833 ( .A(n566), .B(n536), .C(n559), .D(n6172), .E(n537), 
        .F(n557), .Z(n6707) );
  HS65_LS_AOI222X2 U9834 ( .A(n40), .B(n10), .C(n33), .D(n4579), .E(n11), .F(
        n31), .Z(n5114) );
  HS65_LS_AOI222X2 U9835 ( .A(n68), .B(n89), .C(n80), .D(n6356), .E(n70), .F(
        n82), .Z(n6928) );
  HS65_LS_AOI222X2 U9836 ( .A(n247), .B(n268), .C(n259), .D(n4763), .E(n249), 
        .F(n261), .Z(n5336) );
  HS65_LS_AOI222X2 U9837 ( .A(n466), .B(n487), .C(n478), .D(n4802), .E(n468), 
        .F(n480), .Z(n5451) );
  HS65_LS_AOI222X2 U9838 ( .A(n289), .B(n310), .C(n301), .D(n6395), .E(n291), 
        .F(n303), .Z(n7043) );
  HS65_LS_AOI222X2 U9839 ( .A(n493), .B(n522), .C(n515), .D(n6249), .E(n494), 
        .F(n513), .Z(n6812) );
  HS65_LS_AOI222X2 U9840 ( .A(n675), .B(n704), .C(n697), .D(n4656), .E(n676), 
        .F(n695), .Z(n5220) );
  HS65_LS_AOI222X2 U9841 ( .A(n860), .B(n882), .C(n858), .D(n1198), .E(n889), 
        .F(n868), .Z(n1368) );
  HS65_LS_AOI222X2 U9842 ( .A(n778), .B(n800), .C(n776), .D(n1950), .E(n807), 
        .F(n786), .Z(n2120) );
  HS65_LS_AOI222X2 U9843 ( .A(n219), .B(n189), .C(n214), .D(n2963), .E(n190), 
        .F(n212), .Z(n3527) );
  HS65_LS_AOI222X2 U9844 ( .A(n667), .B(n648), .C(n660), .D(n3165), .E(n650), 
        .F(n661), .Z(n3768) );
  HS65_LS_AOI222X2 U9845 ( .A(n589), .B(n619), .C(n608), .D(n593), .E(n616), 
        .F(n601), .Z(n9045) );
  HS65_LS_AOI222X2 U9846 ( .A(n102), .B(n132), .C(n121), .D(n106), .E(n129), 
        .F(n114), .Z(n9103) );
  HS65_LS_AOI222X2 U9847 ( .A(n104), .B(n129), .C(n135), .D(n8194), .E(n105), 
        .F(n137), .Z(n8829) );
  HS65_LS_AOI222X2 U9848 ( .A(n591), .B(n616), .C(n622), .D(n8162), .E(n592), 
        .F(n624), .Z(n8741) );
  HS65_LS_AOI222X2 U9849 ( .A(n443), .B(n424), .C(n436), .D(n3206), .E(n426), 
        .F(n437), .Z(n3885) );
  HS65_LS_AOI222X2 U9850 ( .A(n352), .B(n319), .C(n344), .D(n327), .E(n323), 
        .F(n354), .Z(n8868) );
  HS65_LS_AOI222X2 U9851 ( .A(n393), .B(n369), .C(n401), .D(n8001), .E(n366), 
        .F(n404), .Z(n8306) );
  HS65_LS_AOI222X2 U9852 ( .A(n148), .B(n174), .C(n167), .D(n157), .E(n149), 
        .F(n175), .Z(n3588) );
  HS65_LS_AOI222X2 U9853 ( .A(n920), .B(n901), .C(n926), .D(n904), .E(n918), 
        .F(n910), .Z(n2485) );
  HS65_LS_AOI222X2 U9854 ( .A(n838), .B(n819), .C(n844), .D(n822), .E(n836), 
        .F(n828), .Z(n1733) );
  HS65_LS_AOI222X2 U9855 ( .A(n879), .B(n860), .C(n885), .D(n863), .E(n877), 
        .F(n869), .Z(n1357) );
  HS65_LS_AOI222X2 U9856 ( .A(n797), .B(n778), .C(n803), .D(n781), .E(n795), 
        .F(n787), .Z(n2109) );
  HS65_LSS_XOR2X3 U9857 ( .A(n3544), .B(n452), .Z(n4424) );
  HS65_LSS_XOR2X3 U9858 ( .A(n3219), .B(n275), .Z(n6017) );
  HS65_LS_AOI212X2 U9859 ( .A(n644), .B(n3710), .C(n640), .D(n669), .E(n4289), 
        .Z(n4284) );
  HS65_LS_CB4I6X4 U9860 ( .A(n635), .B(n639), .C(n658), .D(n3782), .Z(n4289)
         );
  HS65_LS_NAND4ABX3 U9861 ( .A(n2419), .B(n2420), .C(n2421), .D(n2422), .Z(
        n2278) );
  HS65_LS_MX41X4 U9862 ( .D0(n918), .S0(n904), .D1(n901), .S1(n921), .D2(n909), 
        .S2(n917), .D3(n929), .S3(n2484), .Z(n2419) );
  HS65_LS_NAND4ABX3 U9863 ( .A(n2480), .B(n2481), .C(n2482), .D(n2483), .Z(
        n2420) );
  HS65_LS_AOI212X2 U9864 ( .A(n899), .B(n2423), .C(n924), .D(n2345), .E(n2424), 
        .Z(n2422) );
  HS65_LS_NAND4ABX3 U9865 ( .A(n1667), .B(n1668), .C(n1669), .D(n1670), .Z(
        n1526) );
  HS65_LS_MX41X4 U9866 ( .D0(n836), .S0(n822), .D1(n819), .S1(n839), .D2(n827), 
        .S2(n835), .D3(n847), .S3(n1732), .Z(n1667) );
  HS65_LS_NAND4ABX3 U9867 ( .A(n1728), .B(n1729), .C(n1730), .D(n1731), .Z(
        n1668) );
  HS65_LS_AOI212X2 U9868 ( .A(n817), .B(n1671), .C(n842), .D(n1593), .E(n1672), 
        .Z(n1670) );
  HS65_LS_NAND4ABX3 U9869 ( .A(n1291), .B(n1292), .C(n1293), .D(n1294), .Z(
        n1150) );
  HS65_LS_NAND4ABX3 U9870 ( .A(n1352), .B(n1353), .C(n1354), .D(n1355), .Z(
        n1292) );
  HS65_LS_MX41X4 U9871 ( .D0(n877), .S0(n863), .D1(n860), .S1(n880), .D2(n868), 
        .S2(n876), .D3(n888), .S3(n1356), .Z(n1291) );
  HS65_LS_AOI212X2 U9872 ( .A(n858), .B(n1295), .C(n883), .D(n1217), .E(n1296), 
        .Z(n1294) );
  HS65_LS_NAND4ABX3 U9873 ( .A(n2043), .B(n2044), .C(n2045), .D(n2046), .Z(
        n1902) );
  HS65_LS_NAND4ABX3 U9874 ( .A(n2104), .B(n2105), .C(n2106), .D(n2107), .Z(
        n2044) );
  HS65_LS_MX41X4 U9875 ( .D0(n795), .S0(n781), .D1(n778), .S1(n798), .D2(n786), 
        .S2(n794), .D3(n806), .S3(n2108), .Z(n2043) );
  HS65_LS_AOI212X2 U9876 ( .A(n776), .B(n2047), .C(n801), .D(n1969), .E(n2048), 
        .Z(n2046) );
  HS65_LSS_XOR2X3 U9877 ( .A(n2813), .B(n7542), .Z(n7615) );
  HS65_LSS_XNOR2X3 U9878 ( .A(n2821), .B(n5950), .Z(n6026) );
  HS65_LSS_XNOR2X3 U9879 ( .A(n2829), .B(n4357), .Z(n4433) );
  HS65_LSS_XOR2X3 U9880 ( .A(n2785), .B(n7542), .Z(n7650) );
  HS65_LS_NAND4ABX3 U9881 ( .A(n4323), .B(n4324), .C(n4325), .D(n4326), .Z(
        n3981) );
  HS65_LS_NOR4ABX2 U9882 ( .A(n4327), .B(n3878), .C(n3398), .D(n3798), .Z(
        n4326) );
  HS65_LS_AOI222X2 U9883 ( .A(n439), .B(n425), .C(n436), .D(n411), .E(n410), 
        .F(n445), .Z(n4325) );
  HS65_LS_NAND4ABX3 U9884 ( .A(n3198), .B(n3838), .C(n3818), .D(n3854), .Z(
        n4323) );
  HS65_LS_NAND4ABX3 U9885 ( .A(n4264), .B(n4265), .C(n4266), .D(n4267), .Z(
        n3960) );
  HS65_LS_AOI222X2 U9886 ( .A(n663), .B(n649), .C(n660), .D(n634), .E(n633), 
        .F(n669), .Z(n4266) );
  HS65_LS_NAND4ABX3 U9887 ( .A(n3157), .B(n3699), .C(n3718), .D(n3737), .Z(
        n4264) );
  HS65_LS_NAND4ABX3 U9888 ( .A(n3344), .B(n3706), .C(n3773), .D(n3321), .Z(
        n4265) );
  HS65_LS_NAND4ABX3 U9889 ( .A(n1814), .B(n1815), .C(n1816), .D(n1817), .Z(
        n1788) );
  HS65_LS_AOI212X2 U9890 ( .A(n817), .B(n1741), .C(n843), .D(n822), .E(n1818), 
        .Z(n1817) );
  HS65_LS_NAND3AX3 U9891 ( .A(n1624), .B(n1711), .C(n1835), .Z(n1815) );
  HS65_LS_MX41X4 U9892 ( .D0(n815), .S0(n844), .D1(n819), .S1(n839), .D2(n836), 
        .S2(n813), .D3(n825), .S3(n837), .Z(n1814) );
  HS65_LS_NAND4ABX3 U9893 ( .A(n2566), .B(n2567), .C(n2568), .D(n2569), .Z(
        n2540) );
  HS65_LS_AOI212X2 U9894 ( .A(n899), .B(n2493), .C(n925), .D(n904), .E(n2570), 
        .Z(n2569) );
  HS65_LS_NAND3AX3 U9895 ( .A(n2376), .B(n2463), .C(n2587), .Z(n2567) );
  HS65_LS_MX41X4 U9896 ( .D0(n897), .S0(n926), .D1(n901), .S1(n921), .D2(n918), 
        .S2(n895), .D3(n907), .S3(n919), .Z(n2566) );
  HS65_LS_NAND4ABX3 U9897 ( .A(n1438), .B(n1439), .C(n1440), .D(n1441), .Z(
        n1412) );
  HS65_LS_NAND3AX3 U9898 ( .A(n1248), .B(n1335), .C(n1459), .Z(n1439) );
  HS65_LS_MX41X4 U9899 ( .D0(n856), .S0(n885), .D1(n860), .S1(n880), .D2(n877), 
        .S2(n854), .D3(n866), .S3(n878), .Z(n1438) );
  HS65_LS_AOI212X2 U9900 ( .A(n858), .B(n1365), .C(n884), .D(n863), .E(n1442), 
        .Z(n1441) );
  HS65_LS_NAND4ABX3 U9901 ( .A(n2190), .B(n2191), .C(n2192), .D(n2193), .Z(
        n2164) );
  HS65_LS_NAND3AX3 U9902 ( .A(n2000), .B(n2087), .C(n2211), .Z(n2191) );
  HS65_LS_MX41X4 U9903 ( .D0(n774), .S0(n803), .D1(n778), .S1(n798), .D2(n795), 
        .S2(n772), .D3(n784), .S3(n796), .Z(n2190) );
  HS65_LS_AOI212X2 U9904 ( .A(n776), .B(n2117), .C(n802), .D(n781), .E(n2194), 
        .Z(n2193) );
  HS65_LS_NAND4ABX3 U9905 ( .A(n4242), .B(n4243), .C(n4244), .D(n4245), .Z(
        n4011) );
  HS65_LS_AOI212X2 U9906 ( .A(n660), .B(n3695), .C(n640), .D(n659), .E(n4246), 
        .Z(n4245) );
  HS65_LS_MX41X4 U9907 ( .D0(n671), .S0(n635), .D1(n667), .S1(n641), .D2(n646), 
        .S2(n662), .D3(n664), .S3(n647), .Z(n4242) );
  HS65_LS_NAND3AX3 U9908 ( .A(n3334), .B(n3751), .C(n4263), .Z(n4243) );
  HS65_LS_NAND4ABX3 U9909 ( .A(n4092), .B(n4093), .C(n4094), .D(n4095), .Z(
        n3996) );
  HS65_LS_NAND3X2 U9910 ( .A(n3266), .B(n3635), .C(n4106), .Z(n4093) );
  HS65_LS_MX41X4 U9911 ( .D0(n177), .S0(n157), .D1(n155), .S1(n174), .D2(n149), 
        .S2(n165), .D3(n172), .S3(n147), .Z(n4092) );
  HS65_LS_AOI212X2 U9912 ( .A(n168), .B(n3596), .C(n156), .D(n167), .E(n4096), 
        .Z(n4095) );
  HS65_LS_NAND4ABX3 U9913 ( .A(n4062), .B(n4063), .C(n4064), .D(n4065), .Z(
        n3934) );
  HS65_LS_AOI212X2 U9914 ( .A(n214), .B(n3451), .C(n201), .D(n213), .E(n4066), 
        .Z(n4065) );
  HS65_LS_MX41X4 U9915 ( .D0(n222), .S0(n202), .D1(n219), .S1(n200), .D2(n194), 
        .S2(n210), .D3(n217), .S3(n192), .Z(n4062) );
  HS65_LS_NAND3AX3 U9916 ( .A(n3107), .B(n3510), .C(n4075), .Z(n4063) );
  HS65_LS_NAND4ABX3 U9917 ( .A(n4301), .B(n4302), .C(n4303), .D(n4304), .Z(
        n4035) );
  HS65_LS_MX41X4 U9918 ( .D0(n447), .S0(n412), .D1(n443), .S1(n417), .D2(n422), 
        .S2(n438), .D3(n440), .S3(n423), .Z(n4301) );
  HS65_LS_NAND3AX3 U9919 ( .A(n3396), .B(n3868), .C(n4322), .Z(n4302) );
  HS65_LS_AOI212X2 U9920 ( .A(n436), .B(n3812), .C(n416), .D(n435), .E(n4305), 
        .Z(n4304) );
  HS65_LS_NOR4ABX2 U9921 ( .A(n4151), .B(n4152), .C(n4153), .D(n4154), .Z(
        n4105) );
  HS65_LS_NAND4ABX3 U9922 ( .A(n3661), .B(n3622), .C(n3607), .D(n2930), .Z(
        n4153) );
  HS65_LS_NAND4ABX3 U9923 ( .A(n3569), .B(n3270), .C(n3595), .D(n3062), .Z(
        n4154) );
  HS65_LS_NOR3AX2 U9924 ( .A(n4159), .B(n3581), .C(n3294), .Z(n4152) );
  HS65_LS_NOR4ABX2 U9925 ( .A(n8961), .B(n8962), .C(n8963), .D(n8964), .Z(
        n8505) );
  HS65_LS_NAND4ABX3 U9926 ( .A(n8027), .B(n8231), .C(n8270), .D(n8121), .Z(
        n8964) );
  HS65_LS_NAND4ABX3 U9927 ( .A(n8103), .B(n8318), .C(n8090), .D(n8965), .Z(
        n8963) );
  HS65_LS_AOI222X2 U9928 ( .A(n403), .B(n369), .C(n378), .D(n398), .E(n377), 
        .F(n404), .Z(n8961) );
  HS65_LS_NOR4ABX2 U9929 ( .A(n4117), .B(n4118), .C(n4119), .D(n4120), .Z(
        n4090) );
  HS65_LS_NAND3AX3 U9930 ( .A(n3260), .B(n3570), .C(n3587), .Z(n4120) );
  HS65_LS_NAND4ABX3 U9931 ( .A(n3659), .B(n3047), .C(n3624), .D(n3649), .Z(
        n4119) );
  HS65_LS_AOI222X2 U9932 ( .A(n143), .B(n180), .C(n160), .D(n166), .E(n158), 
        .F(n174), .Z(n4117) );
  HS65_LS_NOR4ABX2 U9933 ( .A(n2206), .B(n2207), .C(n2208), .D(n2209), .Z(
        n2147) );
  HS65_LS_NAND3AX3 U9934 ( .A(n2099), .B(n1931), .C(n2210), .Z(n2209) );
  HS65_LS_NOR4X4 U9935 ( .A(n1990), .B(n2001), .C(n2009), .D(n2113), .Z(n2207)
         );
  HS65_LS_NAND4ABX3 U9936 ( .A(n1963), .B(n2025), .C(n1944), .D(n2083), .Z(
        n2208) );
  HS65_LS_NOR4ABX2 U9937 ( .A(n1454), .B(n1455), .C(n1456), .D(n1457), .Z(
        n1395) );
  HS65_LS_NAND3AX3 U9938 ( .A(n1347), .B(n1179), .C(n1458), .Z(n1457) );
  HS65_LS_NOR4X4 U9939 ( .A(n1238), .B(n1249), .C(n1257), .D(n1361), .Z(n1455)
         );
  HS65_LS_NAND4ABX3 U9940 ( .A(n1211), .B(n1273), .C(n1192), .D(n1331), .Z(
        n1456) );
  HS65_LS_NOR4ABX2 U9941 ( .A(n1830), .B(n1831), .C(n1832), .D(n1833), .Z(
        n1771) );
  HS65_LS_NAND3AX3 U9942 ( .A(n1723), .B(n1555), .C(n1834), .Z(n1833) );
  HS65_LS_NAND4ABX3 U9943 ( .A(n1587), .B(n1649), .C(n1568), .D(n1707), .Z(
        n1832) );
  HS65_LS_NOR4X4 U9944 ( .A(n1614), .B(n1625), .C(n1633), .D(n1737), .Z(n1831)
         );
  HS65_LS_NOR4ABX2 U9945 ( .A(n2582), .B(n2583), .C(n2584), .D(n2585), .Z(
        n2523) );
  HS65_LS_NAND3AX3 U9946 ( .A(n2475), .B(n2307), .C(n2586), .Z(n2585) );
  HS65_LS_NOR4X4 U9947 ( .A(n2366), .B(n2377), .C(n2385), .D(n2489), .Z(n2583)
         );
  HS65_LS_NAND4ABX3 U9948 ( .A(n2339), .B(n2401), .C(n2320), .D(n2459), .Z(
        n2584) );
  HS65_LSS_XOR2X3 U9949 ( .A(n3010), .B(n7556), .Z(n7559) );
  HS65_LS_NOR4ABX2 U9950 ( .A(n8901), .B(n8902), .C(n8903), .D(n8904), .Z(
        n8879) );
  HS65_LS_NAND4ABX3 U9951 ( .A(n8071), .B(n8620), .C(n8574), .D(n8363), .Z(
        n8904) );
  HS65_LS_NAND4ABX3 U9952 ( .A(n8344), .B(n8534), .C(n8375), .D(n8905), .Z(
        n8903) );
  HS65_LS_AOI222X2 U9953 ( .A(n341), .B(n322), .C(n329), .D(n351), .E(n326), 
        .F(n345), .Z(n8901) );
  HS65_LS_NOR4ABX2 U9954 ( .A(n4283), .B(n4284), .C(n4285), .D(n4286), .Z(
        n2888) );
  HS65_LS_NAND4ABX3 U9955 ( .A(n3160), .B(n3328), .C(n3683), .D(n3746), .Z(
        n4285) );
  HS65_LS_NAND3AX3 U9956 ( .A(n3723), .B(n3765), .C(n3672), .Z(n4286) );
  HS65_LS_AOI222X2 U9957 ( .A(n648), .B(n656), .C(n661), .D(n634), .E(n667), 
        .F(n633), .Z(n4283) );
  HS65_LS_NOR4ABX2 U9958 ( .A(n8889), .B(n8890), .C(n8891), .D(n8892), .Z(
        n7781) );
  HS65_LS_NAND3AX3 U9959 ( .A(n8625), .B(n8606), .C(n8893), .Z(n8892) );
  HS65_LS_MX41X4 U9960 ( .D0(n324), .S0(n358), .D1(n357), .S1(n332), .D2(n341), 
        .S2(n334), .D3(n318), .S3(n351), .Z(n8891) );
  HS65_LS_AOI212X2 U9961 ( .A(n344), .B(n8522), .C(n330), .D(n343), .E(n8894), 
        .Z(n8890) );
  HS65_LS_NOR4ABX2 U9962 ( .A(n8949), .B(n8950), .C(n8951), .D(n8952), .Z(
        n7764) );
  HS65_LS_NAND3X2 U9963 ( .A(n8302), .B(n8239), .C(n8953), .Z(n8952) );
  HS65_LS_MX41X4 U9964 ( .D0(n374), .S0(n395), .D1(n393), .S1(n381), .D2(n403), 
        .S2(n372), .D3(n365), .S3(n398), .Z(n8951) );
  HS65_LS_AOI212X2 U9965 ( .A(n401), .B(n8217), .C(n379), .D(n402), .E(n8954), 
        .Z(n8950) );
  HS65_LS_NOR4ABX2 U9966 ( .A(n8545), .B(n8546), .C(n8547), .D(n8548), .Z(
        n7956) );
  HS65_LS_NAND4ABX3 U9967 ( .A(n8549), .B(n8550), .C(n8551), .D(n8552), .Z(
        n8548) );
  HS65_LS_MX41X4 U9968 ( .D0(n334), .S0(n343), .D1(n357), .S1(n332), .D2(n345), 
        .S2(n319), .D3(n327), .S3(n8553), .Z(n8547) );
  HS65_LS_AOI212X2 U9969 ( .A(n344), .B(n8554), .C(n337), .D(n8333), .E(n8555), 
        .Z(n8546) );
  HS65_LS_NOR4ABX2 U9970 ( .A(n2485), .B(n2486), .C(n2487), .D(n2488), .Z(
        n2294) );
  HS65_LS_NAND4ABX3 U9971 ( .A(n2489), .B(n2490), .C(n2491), .D(n2492), .Z(
        n2488) );
  HS65_LS_MX41X4 U9972 ( .D0(n921), .S0(n908), .D1(n909), .S1(n929), .D2(n907), 
        .S2(n919), .D3(n897), .S3(n916), .Z(n2487) );
  HS65_LS_AOI212X2 U9973 ( .A(n894), .B(n2493), .C(n896), .D(n2494), .E(n2495), 
        .Z(n2486) );
  HS65_LS_NOR4ABX2 U9974 ( .A(n1733), .B(n1734), .C(n1735), .D(n1736), .Z(
        n1542) );
  HS65_LS_NAND4ABX3 U9975 ( .A(n1737), .B(n1738), .C(n1739), .D(n1740), .Z(
        n1736) );
  HS65_LS_MX41X4 U9976 ( .D0(n839), .S0(n826), .D1(n827), .S1(n847), .D2(n825), 
        .S2(n837), .D3(n815), .S3(n834), .Z(n1735) );
  HS65_LS_AOI212X2 U9977 ( .A(n812), .B(n1741), .C(n814), .D(n1742), .E(n1743), 
        .Z(n1734) );
  HS65_LS_NOR4ABX2 U9978 ( .A(n1357), .B(n1358), .C(n1359), .D(n1360), .Z(
        n1166) );
  HS65_LS_NAND4ABX3 U9979 ( .A(n1361), .B(n1362), .C(n1363), .D(n1364), .Z(
        n1360) );
  HS65_LS_MX41X4 U9980 ( .D0(n880), .S0(n867), .D1(n868), .S1(n888), .D2(n866), 
        .S2(n878), .D3(n856), .S3(n875), .Z(n1359) );
  HS65_LS_AOI212X2 U9981 ( .A(n853), .B(n1365), .C(n855), .D(n1366), .E(n1367), 
        .Z(n1358) );
  HS65_LS_NOR4ABX2 U9982 ( .A(n2109), .B(n2110), .C(n2111), .D(n2112), .Z(
        n1918) );
  HS65_LS_NAND4ABX3 U9983 ( .A(n2113), .B(n2114), .C(n2115), .D(n2116), .Z(
        n2112) );
  HS65_LS_MX41X4 U9984 ( .D0(n798), .S0(n785), .D1(n786), .S1(n806), .D2(n784), 
        .S2(n796), .D3(n774), .S3(n793), .Z(n2111) );
  HS65_LS_AOI212X2 U9985 ( .A(n771), .B(n2117), .C(n773), .D(n2118), .E(n2119), 
        .Z(n2110) );
  HS65_LS_NOR4ABX2 U9986 ( .A(n1479), .B(n1480), .C(n1481), .D(n1482), .Z(
        n1123) );
  HS65_LS_NAND4ABX3 U9987 ( .A(n1185), .B(n1242), .C(n1283), .D(n1330), .Z(
        n1481) );
  HS65_LS_AOI222X2 U9988 ( .A(n882), .B(n853), .C(n868), .D(n888), .E(n860), 
        .F(n874), .Z(n1479) );
  HS65_LS_NOR3AX2 U9989 ( .A(n1349), .B(n1272), .C(n1307), .Z(n1480) );
  HS65_LS_NOR4ABX2 U9990 ( .A(n2607), .B(n2608), .C(n2609), .D(n2610), .Z(
        n2251) );
  HS65_LS_NAND4ABX3 U9991 ( .A(n2313), .B(n2370), .C(n2411), .D(n2458), .Z(
        n2609) );
  HS65_LS_AOI222X2 U9992 ( .A(n923), .B(n894), .C(n909), .D(n929), .E(n901), 
        .F(n915), .Z(n2607) );
  HS65_LS_NOR3AX2 U9993 ( .A(n2477), .B(n2400), .C(n2435), .Z(n2608) );
  HS65_LS_NOR4ABX2 U9994 ( .A(n1855), .B(n1856), .C(n1857), .D(n1858), .Z(
        n1499) );
  HS65_LS_NAND4ABX3 U9995 ( .A(n1561), .B(n1618), .C(n1659), .D(n1706), .Z(
        n1857) );
  HS65_LS_AOI222X2 U9996 ( .A(n841), .B(n812), .C(n827), .D(n847), .E(n819), 
        .F(n833), .Z(n1855) );
  HS65_LS_NOR3AX2 U9997 ( .A(n1725), .B(n1648), .C(n1683), .Z(n1856) );
  HS65_LS_NOR4ABX2 U9998 ( .A(n2231), .B(n2232), .C(n2233), .D(n2234), .Z(
        n1875) );
  HS65_LS_NAND4ABX3 U9999 ( .A(n1937), .B(n1994), .C(n2035), .D(n2082), .Z(
        n2233) );
  HS65_LS_AOI222X2 U10000 ( .A(n800), .B(n771), .C(n786), .D(n806), .E(n778), 
        .F(n792), .Z(n2231) );
  HS65_LS_NOR3AX2 U10001 ( .A(n2101), .B(n2024), .C(n2059), .Z(n2232) );
  HS65_LS_NOR4ABX2 U10002 ( .A(n4342), .B(n4343), .C(n4344), .D(n4345), .Z(
        n2843) );
  HS65_LS_NAND4ABX3 U10003 ( .A(n3201), .B(n3390), .C(n3800), .D(n3863), .Z(
        n4344) );
  HS65_LS_AOI222X2 U10004 ( .A(n424), .B(n432), .C(n437), .D(n411), .E(n443), 
        .F(n410), .Z(n4342) );
  HS65_LS_NOR3AX2 U10005 ( .A(n3882), .B(n3789), .C(n3840), .Z(n4343) );
  HS65_LS_NAND4ABX3 U10006 ( .A(n5894), .B(n5895), .C(n5896), .D(n5897), .Z(
        n5556) );
  HS65_LS_AOI222X2 U10007 ( .A(n467), .B(n486), .C(n474), .D(n455), .E(n459), 
        .F(n487), .Z(n5896) );
  HS65_LS_NOR4ABX2 U10008 ( .A(n5477), .B(n4986), .C(n5434), .D(n5410), .Z(
        n5897) );
  HS65_LS_NAND4ABX3 U10009 ( .A(n5371), .B(n5391), .C(n5898), .D(n4998), .Z(
        n5895) );
  HS65_LS_NAND4ABX3 U10010 ( .A(n5835), .B(n5836), .C(n5837), .D(n5838), .Z(
        n5535) );
  HS65_LS_AOI222X2 U10011 ( .A(n248), .B(n267), .C(n255), .D(n236), .E(n240), 
        .F(n268), .Z(n5837) );
  HS65_LS_NOR4ABX2 U10012 ( .A(n5362), .B(n4932), .C(n5319), .D(n5295), .Z(
        n5838) );
  HS65_LS_NAND4ABX3 U10013 ( .A(n5256), .B(n5276), .C(n5839), .D(n4944), .Z(
        n5836) );
  HS65_LS_NAND4ABX3 U10014 ( .A(n5686), .B(n5687), .C(n5688), .D(n5689), .Z(
        n5502) );
  HS65_LS_AOI222X2 U10015 ( .A(n677), .B(n705), .C(n710), .D(n689), .E(n685), 
        .F(n704), .Z(n5688) );
  HS65_LS_NOR4ABX2 U10016 ( .A(n5247), .B(n4856), .C(n5203), .D(n5178), .Z(
        n5689) );
  HS65_LS_NAND4ABX3 U10017 ( .A(n5138), .B(n5159), .C(n5690), .D(n4870), .Z(
        n5687) );
  HS65_LS_NAND4ABX3 U10018 ( .A(n7486), .B(n7487), .C(n7488), .D(n7489), .Z(
        n7148) );
  HS65_LS_AOI222X2 U10019 ( .A(n290), .B(n309), .C(n297), .D(n278), .E(n282), 
        .F(n310), .Z(n7488) );
  HS65_LS_NOR4ABX2 U10020 ( .A(n7069), .B(n6579), .C(n7026), .D(n7002), .Z(
        n7489) );
  HS65_LS_NAND4ABX3 U10021 ( .A(n6963), .B(n6983), .C(n7490), .D(n6591), .Z(
        n7487) );
  HS65_LS_NAND4ABX3 U10022 ( .A(n7427), .B(n7428), .C(n7429), .D(n7430), .Z(
        n7127) );
  HS65_LS_AOI222X2 U10023 ( .A(n69), .B(n88), .C(n76), .D(n57), .E(n61), .F(
        n89), .Z(n7429) );
  HS65_LS_NOR4ABX2 U10024 ( .A(n6954), .B(n6525), .C(n6911), .D(n6887), .Z(
        n7430) );
  HS65_LS_NAND4ABX3 U10025 ( .A(n6848), .B(n6868), .C(n7431), .D(n6537), .Z(
        n7428) );
  HS65_LS_NAND4ABX3 U10026 ( .A(n7278), .B(n7279), .C(n7280), .D(n7281), .Z(
        n7094) );
  HS65_LS_AOI222X2 U10027 ( .A(n495), .B(n523), .C(n528), .D(n507), .E(n503), 
        .F(n522), .Z(n7280) );
  HS65_LS_NOR4ABX2 U10028 ( .A(n6839), .B(n6449), .C(n6795), .D(n6770), .Z(
        n7281) );
  HS65_LS_NAND4ABX3 U10029 ( .A(n6730), .B(n6751), .C(n7282), .D(n6463), .Z(
        n7279) );
  HS65_LS_NAND4ABX3 U10030 ( .A(n5656), .B(n5657), .C(n5658), .D(n5659), .Z(
        n5486) );
  HS65_LS_AOI222X2 U10031 ( .A(n12), .B(n41), .C(n25), .D(n46), .E(n40), .F(
        n21), .Z(n5658) );
  HS65_LS_NOR4ABX2 U10032 ( .A(n5079), .B(n4716), .C(n5056), .D(n5112), .Z(
        n5659) );
  HS65_LS_NAND4ABX3 U10033 ( .A(n5016), .B(n5037), .C(n5660), .D(n4730), .Z(
        n5657) );
  HS65_LS_NAND4ABX3 U10034 ( .A(n7248), .B(n7249), .C(n7250), .D(n7251), .Z(
        n7078) );
  HS65_LS_AOI222X2 U10035 ( .A(n538), .B(n567), .C(n551), .D(n572), .E(n566), 
        .F(n547), .Z(n7250) );
  HS65_LS_NOR4ABX2 U10036 ( .A(n6672), .B(n6309), .C(n6649), .D(n6705), .Z(
        n7251) );
  HS65_LS_NAND4ABX3 U10037 ( .A(n6609), .B(n6630), .C(n7252), .D(n6323), .Z(
        n7249) );
  HS65_LS_NAND4ABX3 U10038 ( .A(n8874), .B(n8875), .C(n8876), .D(n8877), .Z(
        n7783) );
  HS65_LS_NOR4ABX2 U10039 ( .A(n8601), .B(n8587), .C(n8366), .D(n8621), .Z(
        n8877) );
  HS65_LS_AOI222X2 U10040 ( .A(n356), .B(n319), .C(n347), .D(n332), .E(n357), 
        .F(n327), .Z(n8876) );
  HS65_LS_NAND4ABX3 U10041 ( .A(n8517), .B(n8345), .C(n8570), .D(n8878), .Z(
        n8875) );
  HS65_LS_NAND4ABX3 U10042 ( .A(n8500), .B(n8501), .C(n8502), .D(n8503), .Z(
        n7766) );
  HS65_LS_AOI222X2 U10043 ( .A(n394), .B(n367), .C(n387), .D(n381), .E(n393), 
        .F(n375), .Z(n8502) );
  HS65_LS_NOR4ABX2 U10044 ( .A(n8294), .B(n8120), .C(n8287), .D(n8230), .Z(
        n8503) );
  HS65_LS_NAND4ABX3 U10045 ( .A(n8104), .B(n8268), .C(n8212), .D(n8504), .Z(
        n8501) );
  HS65_LS_NAND4ABX3 U10046 ( .A(n8820), .B(n8821), .C(n8822), .D(n8823), .Z(
        n8175) );
  HS65_LS_AOI212X2 U10047 ( .A(n121), .B(n7733), .C(n125), .D(n8824), .E(n8825), .Z(n8823) );
  HS65_LS_AOI222X2 U10048 ( .A(n129), .B(n98), .C(n112), .D(n138), .E(n97), 
        .F(n132), .Z(n8822) );
  HS65_LS_NAND4ABX3 U10049 ( .A(n8826), .B(n8827), .C(n7901), .D(n8828), .Z(
        n8821) );
  HS65_LS_NAND4ABX3 U10050 ( .A(n8732), .B(n8733), .C(n8734), .D(n8735), .Z(
        n8143) );
  HS65_LS_AOI212X2 U10051 ( .A(n608), .B(n7695), .C(n612), .D(n8736), .E(n8737), .Z(n8735) );
  HS65_LS_AOI222X2 U10052 ( .A(n616), .B(n585), .C(n599), .D(n625), .E(n584), 
        .F(n619), .Z(n8734) );
  HS65_LS_NAND4ABX3 U10053 ( .A(n8738), .B(n8739), .C(n7801), .D(n8740), .Z(
        n8733) );
  HS65_LS_NAND4ABX3 U10054 ( .A(n3691), .B(n3692), .C(n3693), .D(n3694), .Z(
        n3140) );
  HS65_LS_NAND4ABX3 U10055 ( .A(n3698), .B(n3699), .C(n3700), .D(n3701), .Z(
        n3692) );
  HS65_LS_AOI222X2 U10056 ( .A(n643), .B(n667), .C(n635), .D(n659), .E(n646), 
        .F(n670), .Z(n3693) );
  HS65_LS_MX41X4 U10057 ( .D0(n641), .S0(n655), .D1(n661), .S1(n634), .D2(n664), .S2(n647), .D3(n671), .S3(n637), .Z(n3691) );
  HS65_LS_NAND4ABX3 U10058 ( .A(n6917), .B(n6918), .C(n6919), .D(n6920), .Z(
        n6331) );
  HS65_LS_AOI212X2 U10059 ( .A(n76), .B(n6921), .C(n86), .D(n6922), .E(n6923), 
        .Z(n6920) );
  HS65_LS_AOI222X2 U10060 ( .A(n89), .B(n63), .C(n60), .D(n79), .E(n66), .F(
        n88), .Z(n6919) );
  HS65_LS_NAND4ABX3 U10061 ( .A(n6924), .B(n6925), .C(n6926), .D(n6927), .Z(
        n6918) );
  HS65_LS_NAND4ABX3 U10062 ( .A(n5325), .B(n5326), .C(n5327), .D(n5328), .Z(
        n4738) );
  HS65_LS_AOI212X2 U10063 ( .A(n255), .B(n5329), .C(n265), .D(n5330), .E(n5331), .Z(n5328) );
  HS65_LS_AOI222X2 U10064 ( .A(n268), .B(n242), .C(n239), .D(n258), .E(n245), 
        .F(n267), .Z(n5327) );
  HS65_LS_NAND4ABX3 U10065 ( .A(n5332), .B(n5333), .C(n5334), .D(n5335), .Z(
        n5326) );
  HS65_LS_NAND4ABX3 U10066 ( .A(n5440), .B(n5441), .C(n5442), .D(n5443), .Z(
        n4777) );
  HS65_LS_AOI212X2 U10067 ( .A(n474), .B(n5444), .C(n484), .D(n5445), .E(n5446), .Z(n5443) );
  HS65_LS_AOI222X2 U10068 ( .A(n487), .B(n461), .C(n458), .D(n477), .E(n464), 
        .F(n486), .Z(n5442) );
  HS65_LS_NAND4ABX3 U10069 ( .A(n5447), .B(n5448), .C(n5449), .D(n5450), .Z(
        n5441) );
  HS65_LS_NAND4ABX3 U10070 ( .A(n7032), .B(n7033), .C(n7034), .D(n7035), .Z(
        n6370) );
  HS65_LS_AOI212X2 U10071 ( .A(n297), .B(n7036), .C(n307), .D(n7037), .E(n7038), .Z(n7035) );
  HS65_LS_AOI222X2 U10072 ( .A(n310), .B(n284), .C(n281), .D(n300), .E(n287), 
        .F(n309), .Z(n7034) );
  HS65_LS_NAND4ABX3 U10073 ( .A(n7039), .B(n7040), .C(n7041), .D(n7042), .Z(
        n7033) );
  HS65_LS_NAND4ABX3 U10074 ( .A(n6801), .B(n6802), .C(n6803), .D(n6804), .Z(
        n6223) );
  HS65_LS_AOI212X2 U10075 ( .A(n528), .B(n6805), .C(n517), .D(n6806), .E(n6807), .Z(n6804) );
  HS65_LS_AOI222X2 U10076 ( .A(n522), .B(n497), .C(n501), .D(n514), .E(n498), 
        .F(n523), .Z(n6803) );
  HS65_LS_NAND4ABX3 U10077 ( .A(n6808), .B(n6809), .C(n6810), .D(n6811), .Z(
        n6802) );
  HS65_LS_NAND4ABX3 U10078 ( .A(n5209), .B(n5210), .C(n5211), .D(n5212), .Z(
        n4630) );
  HS65_LS_AOI212X2 U10079 ( .A(n710), .B(n5213), .C(n699), .D(n5214), .E(n5215), .Z(n5212) );
  HS65_LS_AOI222X2 U10080 ( .A(n704), .B(n679), .C(n683), .D(n696), .E(n680), 
        .F(n705), .Z(n5211) );
  HS65_LS_NAND4ABX3 U10081 ( .A(n5216), .B(n5217), .C(n5218), .D(n5219), .Z(
        n5210) );
  HS65_LS_NAND4ABX3 U10082 ( .A(n3808), .B(n3809), .C(n3810), .D(n3811), .Z(
        n3181) );
  HS65_LS_AOI212X2 U10083 ( .A(n432), .B(n3812), .C(n442), .D(n3813), .E(n3814), .Z(n3811) );
  HS65_LS_NAND4ABX3 U10084 ( .A(n3815), .B(n3816), .C(n3817), .D(n3818), .Z(
        n3809) );
  HS65_LS_MX41X4 U10085 ( .D0(n417), .S0(n431), .D1(n437), .S1(n411), .D2(n440), .S2(n423), .D3(n447), .S3(n414), .Z(n3808) );
  HS65_LS_NAND4ABX3 U10086 ( .A(n3447), .B(n3448), .C(n3449), .D(n3450), .Z(
        n2937) );
  HS65_LS_AOI212X2 U10087 ( .A(n226), .B(n3451), .C(n215), .D(n3452), .E(n3453), .Z(n3450) );
  HS65_LS_AOI222X2 U10088 ( .A(n193), .B(n219), .C(n202), .D(n213), .E(n194), 
        .F(n221), .Z(n3449) );
  HS65_LS_NAND4ABX3 U10089 ( .A(n3455), .B(n3456), .C(n3457), .D(n3458), .Z(
        n3448) );
  HS65_LS_NAND4ABX3 U10090 ( .A(n6680), .B(n6681), .C(n6682), .D(n6683), .Z(
        n6146) );
  HS65_LS_AOI212X2 U10091 ( .A(n572), .B(n6684), .C(n561), .D(n6685), .E(n6686), .Z(n6683) );
  HS65_LS_AOI222X2 U10092 ( .A(n566), .B(n540), .C(n544), .D(n558), .E(n541), 
        .F(n567), .Z(n6682) );
  HS65_LS_NAND4ABX3 U10093 ( .A(n6687), .B(n6688), .C(n6689), .D(n6690), .Z(
        n6681) );
  HS65_LS_NAND4ABX3 U10094 ( .A(n5087), .B(n5088), .C(n5089), .D(n5090), .Z(
        n4553) );
  HS65_LS_AOI212X2 U10095 ( .A(n46), .B(n5091), .C(n35), .D(n5092), .E(n5093), 
        .Z(n5090) );
  HS65_LS_AOI222X2 U10096 ( .A(n40), .B(n14), .C(n18), .D(n32), .E(n15), .F(
        n41), .Z(n5089) );
  HS65_LS_NAND4ABX3 U10097 ( .A(n5094), .B(n5095), .C(n5096), .D(n5097), .Z(
        n5088) );
  HS65_LS_NAND4ABX3 U10098 ( .A(n5722), .B(n5723), .C(n5724), .D(n5725), .Z(
        n5655) );
  HS65_LS_AOI222X2 U10099 ( .A(n10), .B(n46), .C(n21), .D(n31), .E(n40), .F(
        n20), .Z(n5724) );
  HS65_LS_NAND3AX3 U10100 ( .A(n5035), .B(n5078), .C(n5018), .Z(n5723) );
  HS65_LS_NAND4ABX3 U10101 ( .A(n4574), .B(n4717), .C(n5110), .D(n5054), .Z(
        n5722) );
  HS65_LS_NAND4ABX3 U10102 ( .A(n7314), .B(n7315), .C(n7316), .D(n7317), .Z(
        n7247) );
  HS65_LS_AOI222X2 U10103 ( .A(n536), .B(n572), .C(n547), .D(n557), .E(n566), 
        .F(n546), .Z(n7316) );
  HS65_LS_NAND3AX3 U10104 ( .A(n6628), .B(n6671), .C(n6611), .Z(n7315) );
  HS65_LS_NAND4ABX3 U10105 ( .A(n6167), .B(n6310), .C(n6703), .D(n6647), .Z(
        n7314) );
  HS65_LS_NAND4ABX3 U10106 ( .A(n4191), .B(n4192), .C(n4193), .D(n4194), .Z(
        n4061) );
  HS65_LS_NAND4ABX3 U10107 ( .A(n2957), .B(n3441), .C(n3097), .D(n3505), .Z(
        n4191) );
  HS65_LS_AOI222X2 U10108 ( .A(n189), .B(n226), .C(n212), .D(n205), .E(n219), 
        .F(n203), .Z(n4193) );
  HS65_LS_NAND3AX3 U10109 ( .A(n3482), .B(n3428), .C(n3524), .Z(n4192) );
  HS65_LS_NAND4ABX3 U10110 ( .A(n7911), .B(n7912), .C(n7913), .D(n7914), .Z(
        n7728) );
  HS65_LS_NAND4ABX3 U10111 ( .A(n7922), .B(n7923), .C(n7924), .D(n7925), .Z(
        n7911) );
  HS65_LS_AOI222X2 U10112 ( .A(n104), .B(n121), .C(n137), .D(n114), .E(n113), 
        .F(n129), .Z(n7913) );
  HS65_LS_NAND3AX3 U10113 ( .A(n7919), .B(n7920), .C(n7921), .Z(n7912) );
  HS65_LS_NAND4ABX3 U10114 ( .A(n7811), .B(n7812), .C(n7813), .D(n7814), .Z(
        n7690) );
  HS65_LS_NAND4ABX3 U10115 ( .A(n7823), .B(n7824), .C(n7825), .D(n7826), .Z(
        n7811) );
  HS65_LS_AOI222X2 U10116 ( .A(n591), .B(n608), .C(n624), .D(n601), .E(n600), 
        .F(n616), .Z(n7813) );
  HS65_LS_NAND3AX3 U10117 ( .A(n7820), .B(n7821), .C(n7822), .Z(n7812) );
  HS65_LS_NAND4ABX3 U10118 ( .A(n5899), .B(n5900), .C(n5901), .D(n5902), .Z(
        n4507) );
  HS65_LS_AOI222X2 U10119 ( .A(n466), .B(n474), .C(n459), .D(n480), .E(n487), 
        .F(n457), .Z(n5901) );
  HS65_LS_NAND3AX3 U10120 ( .A(n5390), .B(n5432), .C(n5373), .Z(n5900) );
  HS65_LS_NAND4ABX3 U10121 ( .A(n4797), .B(n4987), .C(n5476), .D(n5408), .Z(
        n5899) );
  HS65_LS_NAND4ABX3 U10122 ( .A(n5840), .B(n5841), .C(n5842), .D(n5843), .Z(
        n4461) );
  HS65_LS_AOI222X2 U10123 ( .A(n247), .B(n255), .C(n240), .D(n261), .E(n268), 
        .F(n238), .Z(n5842) );
  HS65_LS_NAND3AX3 U10124 ( .A(n5275), .B(n5317), .C(n5258), .Z(n5841) );
  HS65_LS_NAND4ABX3 U10125 ( .A(n4758), .B(n4933), .C(n5361), .D(n5293), .Z(
        n5840) );
  HS65_LS_NAND4ABX3 U10126 ( .A(n5784), .B(n5785), .C(n5786), .D(n5787), .Z(
        n5685) );
  HS65_LS_AOI222X2 U10127 ( .A(n675), .B(n710), .C(n685), .D(n695), .E(n704), 
        .F(n684), .Z(n5786) );
  HS65_LS_NAND3AX3 U10128 ( .A(n5158), .B(n5201), .C(n5140), .Z(n5785) );
  HS65_LS_NAND4ABX3 U10129 ( .A(n4651), .B(n4857), .C(n5246), .D(n5176), .Z(
        n5784) );
  HS65_LS_NAND4ABX3 U10130 ( .A(n7491), .B(n7492), .C(n7493), .D(n7494), .Z(
        n6100) );
  HS65_LS_AOI222X2 U10131 ( .A(n289), .B(n297), .C(n282), .D(n303), .E(n310), 
        .F(n280), .Z(n7493) );
  HS65_LS_NAND3AX3 U10132 ( .A(n6982), .B(n7024), .C(n6965), .Z(n7492) );
  HS65_LS_NAND4ABX3 U10133 ( .A(n6390), .B(n6580), .C(n7068), .D(n7000), .Z(
        n7491) );
  HS65_LS_NAND4ABX3 U10134 ( .A(n7376), .B(n7377), .C(n7378), .D(n7379), .Z(
        n7277) );
  HS65_LS_AOI222X2 U10135 ( .A(n493), .B(n528), .C(n503), .D(n513), .E(n522), 
        .F(n502), .Z(n7378) );
  HS65_LS_NAND3AX3 U10136 ( .A(n6750), .B(n6793), .C(n6732), .Z(n7377) );
  HS65_LS_NAND4ABX3 U10137 ( .A(n6244), .B(n6450), .C(n6838), .D(n6768), .Z(
        n7376) );
  HS65_LS_NAND4ABX3 U10138 ( .A(n7432), .B(n7433), .C(n7434), .D(n7435), .Z(
        n6054) );
  HS65_LS_AOI222X2 U10139 ( .A(n68), .B(n76), .C(n61), .D(n82), .E(n89), .F(
        n59), .Z(n7434) );
  HS65_LS_NAND3AX3 U10140 ( .A(n6867), .B(n6909), .C(n6850), .Z(n7433) );
  HS65_LS_NAND4ABX3 U10141 ( .A(n6351), .B(n6526), .C(n6953), .D(n6885), .Z(
        n7432) );
  HS65_LS_NAND3X2 U10142 ( .A(n5628), .B(n5629), .C(n5630), .Z(n4508) );
  HS65_LS_NOR3AX2 U10143 ( .A(n4985), .B(n5433), .C(n5418), .Z(n5629) );
  HS65_LS_NOR3X1 U10144 ( .A(n5634), .B(n5397), .C(n5479), .Z(n5628) );
  HS65_LS_AOI212X2 U10145 ( .A(n463), .B(n478), .C(n474), .D(n464), .E(n5631), 
        .Z(n5630) );
  HS65_LS_NAND3X2 U10146 ( .A(n5601), .B(n5602), .C(n5603), .Z(n4462) );
  HS65_LS_NOR3AX2 U10147 ( .A(n4931), .B(n5318), .C(n5303), .Z(n5602) );
  HS65_LS_NOR3X1 U10148 ( .A(n5607), .B(n5282), .C(n5364), .Z(n5601) );
  HS65_LS_AOI212X2 U10149 ( .A(n244), .B(n259), .C(n255), .D(n245), .E(n5604), 
        .Z(n5603) );
  HS65_LS_NAND3X2 U10150 ( .A(n7220), .B(n7221), .C(n7222), .Z(n6101) );
  HS65_LS_NOR3AX2 U10151 ( .A(n6578), .B(n7025), .C(n7010), .Z(n7221) );
  HS65_LS_NOR3X1 U10152 ( .A(n7226), .B(n6989), .C(n7071), .Z(n7220) );
  HS65_LS_AOI212X2 U10153 ( .A(n286), .B(n301), .C(n297), .D(n287), .E(n7223), 
        .Z(n7222) );
  HS65_LS_NAND3X2 U10154 ( .A(n5777), .B(n5778), .C(n5779), .Z(n5579) );
  HS65_LS_NOR3AX2 U10155 ( .A(n4855), .B(n5202), .C(n5187), .Z(n5778) );
  HS65_LS_NOR3X1 U10156 ( .A(n5783), .B(n5165), .C(n5249), .Z(n5777) );
  HS65_LS_AOI212X2 U10157 ( .A(n682), .B(n697), .C(n710), .D(n680), .E(n5780), 
        .Z(n5779) );
  HS65_LS_NAND3X2 U10158 ( .A(n7369), .B(n7370), .C(n7371), .Z(n7171) );
  HS65_LS_NOR3AX2 U10159 ( .A(n6448), .B(n6794), .C(n6779), .Z(n7370) );
  HS65_LS_NOR3X1 U10160 ( .A(n7375), .B(n6757), .C(n6841), .Z(n7369) );
  HS65_LS_AOI212X2 U10161 ( .A(n500), .B(n515), .C(n528), .D(n498), .E(n7372), 
        .Z(n7371) );
  HS65_LS_NAND3X2 U10162 ( .A(n7193), .B(n7194), .C(n7195), .Z(n6055) );
  HS65_LS_NOR3AX2 U10163 ( .A(n6524), .B(n6910), .C(n6895), .Z(n7194) );
  HS65_LS_NOR3X1 U10164 ( .A(n7199), .B(n6874), .C(n6956), .Z(n7193) );
  HS65_LS_AOI212X2 U10165 ( .A(n65), .B(n80), .C(n76), .D(n66), .E(n7196), .Z(
        n7195) );
  HS65_LS_NAND3X2 U10166 ( .A(n4012), .B(n4013), .C(n4014), .Z(n2891) );
  HS65_LS_NOR3AX2 U10167 ( .A(n3326), .B(n3766), .C(n3744), .Z(n4013) );
  HS65_LS_NOR3X1 U10168 ( .A(n4018), .B(n3724), .C(n3686), .Z(n4012) );
  HS65_LS_AOI212X2 U10169 ( .A(n660), .B(n645), .C(n646), .D(n656), .E(n4015), 
        .Z(n4014) );
  HS65_LS_NAND3X2 U10170 ( .A(n4036), .B(n4037), .C(n4038), .Z(n2846) );
  HS65_LS_NOR3X1 U10171 ( .A(n3883), .B(n3389), .C(n3861), .Z(n4037) );
  HS65_LS_NOR3X1 U10172 ( .A(n4042), .B(n3841), .C(n3803), .Z(n4036) );
  HS65_LS_AOI212X2 U10173 ( .A(n436), .B(n421), .C(n422), .D(n432), .E(n4039), 
        .Z(n4038) );
  HS65_LS_NAND3X2 U10174 ( .A(n4184), .B(n4185), .C(n4186), .Z(n3933) );
  HS65_LS_NOR3X1 U10175 ( .A(n3525), .B(n3098), .C(n3503), .Z(n4185) );
  HS65_LS_NOR3X1 U10176 ( .A(n4190), .B(n3481), .C(n3442), .Z(n4184) );
  HS65_LS_AOI212X2 U10177 ( .A(n214), .B(n195), .C(n194), .D(n226), .E(n4187), 
        .Z(n4186) );
  HS65_LS_NAND3X2 U10178 ( .A(n1789), .B(n1790), .C(n1791), .Z(n1502) );
  HS65_LS_NOR3X1 U10179 ( .A(n1726), .B(n1617), .C(n1704), .Z(n1790) );
  HS65_LS_NOR3X1 U10180 ( .A(n1795), .B(n1684), .C(n1662), .Z(n1789) );
  HS65_LS_AOI212X2 U10181 ( .A(n817), .B(n846), .C(n836), .D(n812), .E(n1792), 
        .Z(n1791) );
  HS65_LS_NAND3X2 U10182 ( .A(n2541), .B(n2542), .C(n2543), .Z(n2254) );
  HS65_LS_NOR3X1 U10183 ( .A(n2478), .B(n2369), .C(n2456), .Z(n2542) );
  HS65_LS_NOR3X1 U10184 ( .A(n2547), .B(n2436), .C(n2414), .Z(n2541) );
  HS65_LS_AOI212X2 U10185 ( .A(n899), .B(n928), .C(n918), .D(n894), .E(n2544), 
        .Z(n2543) );
  HS65_LS_NAND3X2 U10186 ( .A(n1413), .B(n1414), .C(n1415), .Z(n1126) );
  HS65_LS_NOR3X1 U10187 ( .A(n1350), .B(n1241), .C(n1328), .Z(n1414) );
  HS65_LS_NOR3X1 U10188 ( .A(n1419), .B(n1308), .C(n1286), .Z(n1413) );
  HS65_LS_AOI212X2 U10189 ( .A(n858), .B(n887), .C(n877), .D(n853), .E(n1416), 
        .Z(n1415) );
  HS65_LS_NAND3X2 U10190 ( .A(n2165), .B(n2166), .C(n2167), .Z(n1878) );
  HS65_LS_NOR3X1 U10191 ( .A(n2102), .B(n1993), .C(n2080), .Z(n2166) );
  HS65_LS_NOR3X1 U10192 ( .A(n2171), .B(n2060), .C(n2038), .Z(n2165) );
  HS65_LS_AOI212X2 U10193 ( .A(n776), .B(n805), .C(n795), .D(n771), .E(n2168), 
        .Z(n2167) );
  HS65_LS_NAND3X2 U10194 ( .A(n8971), .B(n8972), .C(n8973), .Z(n8651) );
  HS65_LS_NOR3X1 U10195 ( .A(n8304), .B(n8117), .C(n8281), .Z(n8972) );
  HS65_LS_NOR3AX2 U10196 ( .A(n8240), .B(n8979), .C(n8263), .Z(n8971) );
  HS65_LS_AOI212X2 U10197 ( .A(n401), .B(n373), .C(n372), .D(n387), .E(n8974), 
        .Z(n8973) );
  HS65_LS_NAND3X2 U10198 ( .A(n7926), .B(n7927), .C(n7928), .Z(n7658) );
  HS65_LS_NOR3AX2 U10199 ( .A(n7934), .B(n7935), .C(n7936), .Z(n7927) );
  HS65_LS_NOR3AX2 U10200 ( .A(n7937), .B(n7938), .C(n7939), .Z(n7926) );
  HS65_LS_AOI212X2 U10201 ( .A(n135), .B(n99), .C(n121), .D(n97), .E(n7929), 
        .Z(n7928) );
  HS65_LS_NAND3X2 U10202 ( .A(n7827), .B(n7828), .C(n7829), .Z(n7630) );
  HS65_LS_NOR3AX2 U10203 ( .A(n7835), .B(n7836), .C(n7837), .Z(n7828) );
  HS65_LS_NOR3AX2 U10204 ( .A(n7838), .B(n7839), .C(n7840), .Z(n7827) );
  HS65_LS_AOI212X2 U10205 ( .A(n622), .B(n586), .C(n608), .D(n584), .E(n7830), 
        .Z(n7829) );
  HS65_LS_NAND4ABX3 U10206 ( .A(n8518), .B(n8519), .C(n8520), .D(n8521), .Z(
        n8054) );
  HS65_LS_AOI212X2 U10207 ( .A(n347), .B(n8522), .C(n350), .D(n8523), .E(n8524), .Z(n8521) );
  HS65_LS_AOI222X2 U10208 ( .A(n335), .B(n357), .C(n324), .D(n343), .E(n356), 
        .F(n334), .Z(n8520) );
  HS65_LS_NAND4ABX3 U10209 ( .A(n8526), .B(n8527), .C(n8528), .D(n8529), .Z(
        n8519) );
  HS65_LS_IVX2 U10210 ( .A(n2893), .Z(n639) );
  HS65_LS_NAND4ABX3 U10211 ( .A(n7767), .B(n7768), .C(n7769), .D(n7770), .Z(
        n2908) );
  HS65_LS_MX41X4 U10212 ( .D0(n318), .S0(n352), .D1(n343), .S1(n322), .D2(n335), .S2(n349), .D3(n323), .S3(n344), .Z(n7767) );
  HS65_LS_NOR4ABX2 U10213 ( .A(n7771), .B(n7772), .C(n7773), .D(n7774), .Z(
        n7770) );
  HS65_LS_MX41X4 U10214 ( .D0(n351), .S0(n337), .D1(n331), .S1(n346), .D2(n329), .S2(n353), .D3(n336), .S3(n7784), .Z(n7768) );
  HS65_LS_IVX2 U10215 ( .A(n3015), .Z(n317) );
  HS65_LS_NAND4ABX3 U10216 ( .A(n8213), .B(n8214), .C(n8215), .D(n8216), .Z(
        n8012) );
  HS65_LS_AOI212X2 U10217 ( .A(n387), .B(n8217), .C(n397), .D(n8218), .E(n8219), .Z(n8216) );
  HS65_LS_AOI222X2 U10218 ( .A(n370), .B(n393), .C(n374), .D(n402), .E(n394), 
        .F(n372), .Z(n8215) );
  HS65_LS_MX41X4 U10219 ( .D0(n381), .S0(n386), .D1(n375), .S1(n404), .D2(n365), .S2(n398), .D3(n395), .S3(n380), .Z(n8213) );
  HS65_LS_NOR2X2 U10220 ( .A(n179), .B(n172), .Z(n3051) );
  HS65_LSS_XOR2X3 U10221 ( .A(n3222), .B(n451), .Z(n4373) );
  HS65_LSS_XOR2X3 U10222 ( .A(n3018), .B(n274), .Z(n5966) );
  HS65_LS_NAND4ABX3 U10223 ( .A(n6851), .B(n6852), .C(n6853), .D(n6854), .Z(
        n6193) );
  HS65_LS_NAND4ABX3 U10224 ( .A(n6912), .B(n6913), .C(n6914), .D(n6915), .Z(
        n6852) );
  HS65_LS_MX41X4 U10225 ( .D0(n66), .S0(n79), .D1(n57), .S1(n89), .D2(n69), 
        .S2(n82), .D3(n61), .S3(n6916), .Z(n6851) );
  HS65_LS_AOI212X2 U10226 ( .A(n80), .B(n6855), .C(n64), .D(n6489), .E(n6856), 
        .Z(n6854) );
  HS65_LS_NAND4ABX3 U10227 ( .A(n5259), .B(n5260), .C(n5261), .D(n5262), .Z(
        n4600) );
  HS65_LS_NAND4ABX3 U10228 ( .A(n5320), .B(n5321), .C(n5322), .D(n5323), .Z(
        n5260) );
  HS65_LS_MX41X4 U10229 ( .D0(n245), .S0(n258), .D1(n236), .S1(n268), .D2(n248), .S2(n261), .D3(n240), .S3(n5324), .Z(n5259) );
  HS65_LS_AOI212X2 U10230 ( .A(n259), .B(n5263), .C(n243), .D(n4896), .E(n5264), .Z(n5262) );
  HS65_LS_NAND4ABX3 U10231 ( .A(n5374), .B(n5375), .C(n5376), .D(n5377), .Z(
        n4612) );
  HS65_LS_NAND4ABX3 U10232 ( .A(n5435), .B(n5436), .C(n5437), .D(n5438), .Z(
        n5375) );
  HS65_LS_MX41X4 U10233 ( .D0(n464), .S0(n477), .D1(n455), .S1(n487), .D2(n467), .S2(n480), .D3(n459), .S3(n5439), .Z(n5374) );
  HS65_LS_AOI212X2 U10234 ( .A(n478), .B(n5378), .C(n462), .D(n4950), .E(n5379), .Z(n5377) );
  HS65_LS_NAND4ABX3 U10235 ( .A(n6966), .B(n6967), .C(n6968), .D(n6969), .Z(
        n6205) );
  HS65_LS_NAND4ABX3 U10236 ( .A(n7027), .B(n7028), .C(n7029), .D(n7030), .Z(
        n6967) );
  HS65_LS_MX41X4 U10237 ( .D0(n287), .S0(n300), .D1(n278), .S1(n310), .D2(n290), .S2(n303), .D3(n282), .S3(n7031), .Z(n6966) );
  HS65_LS_AOI212X2 U10238 ( .A(n301), .B(n6970), .C(n285), .D(n6543), .E(n6971), .Z(n6969) );
  HS65_LS_NAND4ABX3 U10239 ( .A(n5141), .B(n5142), .C(n5143), .D(n5144), .Z(
        n4542) );
  HS65_LS_NAND4ABX3 U10240 ( .A(n5204), .B(n5205), .C(n5206), .D(n5207), .Z(
        n5142) );
  HS65_LS_MX41X4 U10241 ( .D0(n680), .S0(n696), .D1(n689), .S1(n704), .D2(n677), .S2(n695), .D3(n685), .S3(n5208), .Z(n5141) );
  HS65_LS_AOI212X2 U10242 ( .A(n697), .B(n5145), .C(n681), .D(n4818), .E(n5146), .Z(n5144) );
  HS65_LS_NAND4ABX3 U10243 ( .A(n6733), .B(n6734), .C(n6735), .D(n6736), .Z(
        n6135) );
  HS65_LS_NAND4ABX3 U10244 ( .A(n6796), .B(n6797), .C(n6798), .D(n6799), .Z(
        n6734) );
  HS65_LS_MX41X4 U10245 ( .D0(n498), .S0(n514), .D1(n507), .S1(n522), .D2(n495), .S2(n513), .D3(n503), .S3(n6800), .Z(n6733) );
  HS65_LS_AOI212X2 U10246 ( .A(n515), .B(n6737), .C(n499), .D(n6411), .E(n6738), .Z(n6736) );
  HS65_LS_NAND4ABX3 U10247 ( .A(n6612), .B(n6613), .C(n6614), .D(n6615), .Z(
        n6079) );
  HS65_LS_NAND4ABX3 U10248 ( .A(n6675), .B(n6676), .C(n6677), .D(n6678), .Z(
        n6613) );
  HS65_LS_MX41X4 U10249 ( .D0(n541), .S0(n558), .D1(n566), .S1(n551), .D2(n538), .S2(n557), .D3(n547), .S3(n6679), .Z(n6612) );
  HS65_LS_AOI212X2 U10250 ( .A(n559), .B(n6616), .C(n542), .D(n6271), .E(n6617), .Z(n6615) );
  HS65_LS_NAND4ABX3 U10251 ( .A(n5019), .B(n5020), .C(n5021), .D(n5022), .Z(
        n4486) );
  HS65_LS_NAND4ABX3 U10252 ( .A(n5082), .B(n5083), .C(n5084), .D(n5085), .Z(
        n5020) );
  HS65_LS_MX41X4 U10253 ( .D0(n15), .S0(n32), .D1(n40), .S1(n25), .D2(n12), 
        .S2(n31), .D3(n21), .S3(n5086), .Z(n5019) );
  HS65_LS_AOI212X2 U10254 ( .A(n33), .B(n5023), .C(n16), .D(n4678), .E(n5024), 
        .Z(n5022) );
  HS65_LS_NAND4ABX3 U10255 ( .A(n8684), .B(n8685), .C(n8686), .D(n8687), .Z(
        n7975) );
  HS65_LS_NAND4ABX3 U10256 ( .A(n8729), .B(n8730), .C(n8731), .D(n7807), .Z(
        n8685) );
  HS65_LS_AOI212X2 U10257 ( .A(n622), .B(n8688), .C(n583), .D(n8388), .E(n8689), .Z(n8687) );
  HS65_LS_MX41X4 U10258 ( .D0(n584), .S0(n625), .D1(n593), .S1(n616), .D2(n589), .S2(n624), .D3(n601), .S3(n7815), .Z(n8684) );
  HS65_LS_NAND4ABX3 U10259 ( .A(n8772), .B(n8773), .C(n8774), .D(n8775), .Z(
        n7988) );
  HS65_LS_NAND4ABX3 U10260 ( .A(n8817), .B(n8818), .C(n8819), .D(n7907), .Z(
        n8773) );
  HS65_LS_AOI212X2 U10261 ( .A(n135), .B(n8776), .C(n96), .D(n8448), .E(n8777), 
        .Z(n8775) );
  HS65_LS_MX41X4 U10262 ( .D0(n97), .S0(n138), .D1(n106), .S1(n129), .D2(n102), 
        .S2(n137), .D3(n114), .S3(n7915), .Z(n8772) );
  HS65_LS_NAND2X2 U10263 ( .A(n350), .B(n319), .Z(n8065) );
  HS65_LS_NOR2X2 U10264 ( .A(n170), .B(n165), .Z(n2929) );
  HS65_LS_NOR2X2 U10265 ( .A(n826), .B(n817), .Z(n1753) );
  HS65_LS_NOR2X2 U10266 ( .A(n908), .B(n899), .Z(n2505) );
  HS65_LS_NOR2X2 U10267 ( .A(n701), .B(n693), .Z(n4545) );
  HS65_LS_NOR2X2 U10268 ( .A(n483), .B(n479), .Z(n4614) );
  HS65_LS_NOR2X2 U10269 ( .A(n306), .B(n302), .Z(n6207) );
  HS65_LS_NOR2X2 U10270 ( .A(n85), .B(n81), .Z(n6195) );
  HS65_LS_NOR2X2 U10271 ( .A(n519), .B(n511), .Z(n6138) );
  HS65_LS_NOR2X2 U10272 ( .A(n264), .B(n260), .Z(n4602) );
  HS65_LS_NOR2X2 U10273 ( .A(n867), .B(n858), .Z(n1377) );
  HS65_LS_NOR2X2 U10274 ( .A(n785), .B(n776), .Z(n2129) );
  HS65_LS_NOR3AX2 U10275 ( .A(n2889), .B(n2890), .C(n2891), .Z(n2883) );
  HS65_LS_NOR3AX2 U10276 ( .A(n2844), .B(n2845), .C(n2846), .Z(n2838) );
  HS65_LS_NOR3AX2 U10277 ( .A(n3910), .B(n4061), .C(n3933), .Z(n4176) );
  HS65_LS_NOR2X2 U10278 ( .A(n563), .B(n555), .Z(n6082) );
  HS65_LS_NOR2X2 U10279 ( .A(n37), .B(n29), .Z(n4489) );
  HS65_LS_NOR2X2 U10280 ( .A(n182), .B(n168), .Z(n3586) );
  HS65_LS_NOR2X2 U10281 ( .A(n441), .B(n438), .Z(n3008) );
  HS65_LS_NOR2X2 U10282 ( .A(n614), .B(n623), .Z(n7641) );
  HS65_LS_NOR2X2 U10283 ( .A(n396), .B(n403), .Z(n7863) );
  HS65_LS_NOR2X2 U10284 ( .A(n665), .B(n662), .Z(n2990) );
  HS65_LS_NOR2X2 U10285 ( .A(n216), .B(n210), .Z(n2879) );
  HS65_LS_NOR2X2 U10286 ( .A(n431), .B(n436), .Z(n3894) );
  HS65_LS_NOR2X2 U10287 ( .A(n228), .B(n214), .Z(n3537) );
  HS65_LS_OAI13X1 U10288 ( .A(n897), .B(n900), .C(n899), .D(n917), .Z(n2352)
         );
  HS65_LS_OAI13X1 U10289 ( .A(n815), .B(n818), .C(n817), .D(n835), .Z(n1600)
         );
  HS65_LS_NOR2X2 U10290 ( .A(n346), .B(n344), .Z(n8543) );
  HS65_LS_NOR2X2 U10291 ( .A(n353), .B(n341), .Z(n7965) );
  HS65_LS_NOR3AX2 U10292 ( .A(n8082), .B(n8013), .C(n7867), .Z(n8076) );
  HS65_LS_NOR2X2 U10293 ( .A(n386), .B(n401), .Z(n8316) );
  HS65_LS_OAI13X1 U10294 ( .A(n856), .B(n859), .C(n858), .D(n876), .Z(n1224)
         );
  HS65_LS_OAI13X1 U10295 ( .A(n774), .B(n777), .C(n776), .D(n794), .Z(n1976)
         );
  HS65_LS_NOR2X2 U10296 ( .A(n655), .B(n660), .Z(n3777) );
  HS65_LS_NAND4ABX3 U10297 ( .A(n8083), .B(n8084), .C(n8085), .D(n8086), .Z(
        n7867) );
  HS65_LS_NOR3AX2 U10298 ( .A(n8087), .B(n8088), .C(n8089), .Z(n8086) );
  HS65_LS_AOI222X2 U10299 ( .A(n370), .B(n396), .C(n393), .D(n372), .E(n371), 
        .F(n388), .Z(n8085) );
  HS65_LS_NAND3X2 U10300 ( .A(n8090), .B(n8091), .C(n8092), .Z(n8084) );
  HS65_LS_OAI13X1 U10301 ( .A(n614), .B(n620), .C(n622), .D(n589), .Z(n8396)
         );
  HS65_LS_OAI13X1 U10302 ( .A(n127), .B(n133), .C(n135), .D(n102), .Z(n8456)
         );
  HS65_LS_NAND4ABX3 U10303 ( .A(n8530), .B(n8531), .C(n8532), .D(n8533), .Z(
        n8337) );
  HS65_LS_NOR3X1 U10304 ( .A(n8534), .B(n8535), .C(n8536), .Z(n8533) );
  HS65_LS_AOI222X2 U10305 ( .A(n357), .B(n322), .C(n344), .D(n8043), .E(n321), 
        .F(n345), .Z(n8532) );
  HS65_LS_NAND4ABX3 U10306 ( .A(n8537), .B(n8538), .C(n8539), .D(n8540), .Z(
        n8531) );
  HS65_LS_OAI13X1 U10307 ( .A(n447), .B(n441), .C(n436), .D(n425), .Z(n3372)
         );
  HS65_LS_OAI13X1 U10308 ( .A(n222), .B(n216), .C(n214), .D(n191), .Z(n3081)
         );
  HS65_LS_OAI13X1 U10309 ( .A(n43), .B(n33), .C(n37), .D(n12), .Z(n4701) );
  HS65_LS_OAI13X1 U10310 ( .A(n569), .B(n559), .C(n563), .D(n538), .Z(n6294)
         );
  HS65_LS_OAI13X1 U10311 ( .A(n87), .B(n80), .C(n85), .D(n69), .Z(n6510) );
  HS65_LS_OAI13X1 U10312 ( .A(n308), .B(n301), .C(n306), .D(n290), .Z(n6564)
         );
  HS65_LS_OAI13X1 U10313 ( .A(n485), .B(n478), .C(n483), .D(n467), .Z(n4971)
         );
  HS65_LS_OAI13X1 U10314 ( .A(n266), .B(n259), .C(n264), .D(n248), .Z(n4917)
         );
  HS65_LS_OAI13X1 U10315 ( .A(n707), .B(n697), .C(n701), .D(n677), .Z(n4841)
         );
  HS65_LS_OAI13X1 U10316 ( .A(n525), .B(n515), .C(n519), .D(n495), .Z(n6434)
         );
  HS65_LS_OAI13X1 U10317 ( .A(n358), .B(n353), .C(n344), .D(n319), .Z(n8342)
         );
  HS65_LS_OAI13X1 U10318 ( .A(n395), .B(n396), .C(n401), .D(n367), .Z(n8101)
         );
  HS65_LS_NAND4ABX3 U10319 ( .A(n4069), .B(n4070), .C(n4071), .D(n4072), .Z(
        n3908) );
  HS65_LS_NAND4ABX3 U10320 ( .A(n3119), .B(n3083), .C(n2956), .D(n3096), .Z(
        n4070) );
  HS65_LS_NOR4ABX2 U10321 ( .A(n3516), .B(n3471), .C(n3487), .D(n3507), .Z(
        n4072) );
  HS65_LS_NAND4ABX3 U10322 ( .A(n3540), .B(n3453), .C(n4073), .D(n3439), .Z(
        n4069) );
  HS65_LS_OAI13X1 U10323 ( .A(n671), .B(n665), .C(n660), .D(n649), .Z(n3310)
         );
  HS65_LS_NAND4ABX3 U10324 ( .A(n3573), .B(n3574), .C(n3575), .D(n3576), .Z(
        n3238) );
  HS65_LS_NOR3X1 U10325 ( .A(n3577), .B(n3578), .C(n3579), .Z(n3576) );
  HS65_LS_NAND4ABX3 U10326 ( .A(n3580), .B(n3581), .C(n3582), .D(n3583), .Z(
        n3574) );
  HS65_LS_AOI222X2 U10327 ( .A(n143), .B(n174), .C(n168), .D(n3055), .E(n166), 
        .F(n144), .Z(n3575) );
  HS65_LS_OAI13X1 U10328 ( .A(n177), .B(n168), .C(n170), .D(n145), .Z(n3243)
         );
  HS65_LS_IVX2 U10329 ( .A(n2807), .Z(n232) );
  HS65_LS_IVX2 U10330 ( .A(n2799), .Z(n52) );
  HS65_LS_NAND2X2 U10331 ( .A(n378), .B(n386), .Z(n8212) );
  HS65_LS_NOR3AX2 U10332 ( .A(n7973), .B(n8143), .C(n8144), .Z(n8139) );
  HS65_LS_NOR3AX2 U10333 ( .A(n7986), .B(n8175), .C(n8176), .Z(n8171) );
  HS65_LS_NOR3AX2 U10334 ( .A(n8391), .B(n7972), .C(n8144), .Z(n8386) );
  HS65_LS_NOR3AX2 U10335 ( .A(n4484), .B(n4553), .C(n4554), .Z(n4549) );
  HS65_LS_NOR3AX2 U10336 ( .A(n6077), .B(n6146), .C(n6147), .Z(n6142) );
  HS65_LS_NOR3AX2 U10337 ( .A(n6191), .B(n6331), .C(n6332), .Z(n6327) );
  HS65_LS_NOR3AX2 U10338 ( .A(n4610), .B(n4777), .C(n4778), .Z(n4773) );
  HS65_LS_NOR3AX2 U10339 ( .A(n6203), .B(n6370), .C(n6371), .Z(n6366) );
  HS65_LS_NOR3AX2 U10340 ( .A(n4598), .B(n4738), .C(n4739), .Z(n4734) );
  HS65_LS_NOR3AX2 U10341 ( .A(n4540), .B(n4630), .C(n4631), .Z(n4626) );
  HS65_LS_NOR3AX2 U10342 ( .A(n6133), .B(n6223), .C(n6224), .Z(n6219) );
  HS65_LS_NOR3AX2 U10343 ( .A(n7706), .B(n7707), .C(n7708), .Z(n7705) );
  HS65_LS_NOR3AX2 U10344 ( .A(n7744), .B(n7745), .C(n7746), .Z(n7743) );
  HS65_LS_NOR3AX2 U10345 ( .A(n4705), .B(n4482), .C(n4706), .Z(n4699) );
  HS65_LS_NOR3AX2 U10346 ( .A(n6298), .B(n6075), .C(n6299), .Z(n6292) );
  HS65_LS_NOR3AX2 U10347 ( .A(n2996), .B(n3181), .C(n3182), .Z(n3177) );
  HS65_LS_NOR3AX2 U10348 ( .A(n3367), .B(n2999), .C(n3182), .Z(n3362) );
  HS65_LS_NOR3AX2 U10349 ( .A(n6514), .B(n6189), .C(n6515), .Z(n6508) );
  HS65_LS_NOR3AX2 U10350 ( .A(n6568), .B(n6201), .C(n6569), .Z(n6562) );
  HS65_LS_NOR3AX2 U10351 ( .A(n4975), .B(n4608), .C(n4976), .Z(n4969) );
  HS65_LS_NOR3AX2 U10352 ( .A(n4921), .B(n4596), .C(n4922), .Z(n4915) );
  HS65_LS_NOR3AX2 U10353 ( .A(n4845), .B(n4538), .C(n4846), .Z(n4839) );
  HS65_LS_NOR3AX2 U10354 ( .A(n6438), .B(n6131), .C(n6439), .Z(n6432) );
  HS65_LS_NOR3AX2 U10355 ( .A(n3305), .B(n2981), .C(n3141), .Z(n3300) );
  HS65_LS_NOR3AX2 U10356 ( .A(n2978), .B(n3140), .C(n3141), .Z(n3136) );
  HS65_LS_NOR3AX2 U10357 ( .A(n2866), .B(n2937), .C(n2938), .Z(n2933) );
  HS65_LS_NOR3AX2 U10358 ( .A(n3076), .B(n2869), .C(n2938), .Z(n3070) );
  HS65_LS_NOR3AX2 U10359 ( .A(n8347), .B(n7951), .C(n8348), .Z(n8340) );
  HS65_LS_NOR3AX2 U10360 ( .A(n2916), .B(n3238), .C(n3030), .Z(n3232) );
  HS65_LS_NOR3AX2 U10361 ( .A(n3490), .B(n2954), .C(n3526), .Z(n4075) );
  HS65_LS_NOR3AX2 U10362 ( .A(n7699), .B(n7700), .C(n7701), .Z(n7693) );
  HS65_LS_AO12X4 U10363 ( .A(n611), .B(n583), .C(n7702), .Z(n7700) );
  HS65_LS_NOR3AX2 U10364 ( .A(n7737), .B(n7738), .C(n7739), .Z(n7731) );
  HS65_LS_AO12X4 U10365 ( .A(n124), .B(n96), .C(n7740), .Z(n7738) );
  HS65_LS_NOR3X1 U10366 ( .A(n7810), .B(n7630), .C(n7690), .Z(n7790) );
  HS65_LS_IVX2 U10367 ( .A(n7964), .Z(n329) );
  HS65_LS_NOR3X1 U10368 ( .A(n4506), .B(n4507), .C(n4508), .Z(n4500) );
  HS65_LS_NOR3X1 U10369 ( .A(n4460), .B(n4461), .C(n4462), .Z(n4454) );
  HS65_LS_NOR3X1 U10370 ( .A(n6099), .B(n6100), .C(n6101), .Z(n6093) );
  HS65_LS_NOR3X1 U10371 ( .A(n5503), .B(n5685), .C(n5579), .Z(n5769) );
  HS65_LS_NOR3X1 U10372 ( .A(n7095), .B(n7277), .C(n7171), .Z(n7361) );
  HS65_LS_NOR3X1 U10373 ( .A(n6053), .B(n6054), .C(n6055), .Z(n6047) );
  HS65_LS_NOR3X1 U10374 ( .A(n5487), .B(n5655), .C(n5514), .Z(n5707) );
  HS65_LS_NOR3X1 U10375 ( .A(n7079), .B(n7247), .C(n7106), .Z(n7299) );
  HS65_LS_NOR3X1 U10376 ( .A(n7782), .B(n8632), .C(n8633), .Z(n8628) );
  HS65_LSS_XOR2X3 U10377 ( .A(n3220), .B(n451), .Z(n4384) );
  HS65_LSS_XOR2X3 U10378 ( .A(n3016), .B(n274), .Z(n5977) );
  HS65_LS_NOR3X1 U10379 ( .A(n1124), .B(n1125), .C(n1126), .Z(n1118) );
  HS65_LS_NOR3X1 U10380 ( .A(n1500), .B(n1501), .C(n1502), .Z(n1494) );
  HS65_LS_NOR3X1 U10381 ( .A(n2252), .B(n2253), .C(n2254), .Z(n2246) );
  HS65_LS_NOR3X1 U10382 ( .A(n1876), .B(n1877), .C(n1878), .Z(n1870) );
  HS65_LS_NOR3X1 U10383 ( .A(n7765), .B(n8499), .C(n8651), .Z(n8647) );
  HS65_LS_NOR3X1 U10384 ( .A(n3927), .B(n4098), .C(n3995), .Z(n4114) );
  HS65_LS_NOR3AX2 U10385 ( .A(n6546), .B(n6371), .C(n6202), .Z(n6541) );
  HS65_LS_NOR3AX2 U10386 ( .A(n4953), .B(n4778), .C(n4609), .Z(n4948) );
  HS65_LS_NOR3AX2 U10387 ( .A(n4822), .B(n4631), .C(n4539), .Z(n4816) );
  HS65_LS_NOR3AX2 U10388 ( .A(n6415), .B(n6224), .C(n6132), .Z(n6409) );
  HS65_LS_NOR3AX2 U10389 ( .A(n3732), .B(n3156), .C(n3767), .Z(n4263) );
  HS65_LS_NOR4ABX2 U10390 ( .A(n7302), .B(n7303), .C(n7304), .D(n7305), .Z(
        n7259) );
  HS65_LS_NAND4ABX3 U10391 ( .A(n6322), .B(n6627), .C(n6159), .D(n6690), .Z(
        n7305) );
  HS65_LS_NAND4ABX3 U10392 ( .A(n6701), .B(n6282), .C(n7306), .D(n6717), .Z(
        n7304) );
  HS65_LS_AOI222X2 U10393 ( .A(n538), .B(n572), .C(n551), .D(n569), .E(n537), 
        .F(n574), .Z(n7302) );
  HS65_LS_NOR4ABX2 U10394 ( .A(n5710), .B(n5711), .C(n5712), .D(n5713), .Z(
        n5667) );
  HS65_LS_NAND4ABX3 U10395 ( .A(n4729), .B(n5034), .C(n4566), .D(n5097), .Z(
        n5713) );
  HS65_LS_NAND4ABX3 U10396 ( .A(n5108), .B(n4689), .C(n5714), .D(n5124), .Z(
        n5712) );
  HS65_LS_AOI222X2 U10397 ( .A(n12), .B(n46), .C(n25), .D(n43), .E(n11), .F(
        n48), .Z(n5710) );
  HS65_LS_NOR4ABX2 U10398 ( .A(n8906), .B(n8907), .C(n8908), .D(n8909), .Z(
        n8631) );
  HS65_LS_NAND4ABX3 U10399 ( .A(n8368), .B(n8072), .C(n8566), .D(n8529), .Z(
        n8909) );
  HS65_LS_NAND4ABX3 U10400 ( .A(n8624), .B(n8535), .C(n8376), .D(n8910), .Z(
        n8908) );
  HS65_LS_AOI222X2 U10401 ( .A(n347), .B(n319), .C(n358), .D(n332), .E(n321), 
        .F(n346), .Z(n8906) );
  HS65_LS_NOR4ABX2 U10402 ( .A(n8966), .B(n8967), .C(n8968), .D(n8969), .Z(
        n8650) );
  HS65_LS_NAND4ABX3 U10403 ( .A(n8126), .B(n8029), .C(n8262), .D(n8224), .Z(
        n8969) );
  HS65_LS_NAND4ABX3 U10404 ( .A(n8237), .B(n8320), .C(n8091), .D(n8970), .Z(
        n8968) );
  HS65_LS_AOI222X2 U10405 ( .A(n387), .B(n367), .C(n395), .D(n381), .E(n366), 
        .F(n386), .Z(n8966) );
  HS65_LS_NOR4ABX2 U10406 ( .A(n4179), .B(n4180), .C(n4181), .D(n4182), .Z(
        n4067) );
  HS65_LS_NAND4ABX3 U10407 ( .A(n3480), .B(n2958), .C(n3110), .D(n3457), .Z(
        n4182) );
  HS65_LS_NAND4ABX3 U10408 ( .A(n4183), .B(n3542), .C(n3440), .D(n3120), .Z(
        n4181) );
  HS65_LS_AOI222X2 U10409 ( .A(n191), .B(n226), .C(n222), .D(n200), .E(n190), 
        .F(n228), .Z(n4179) );
  HS65_LS_NAND4ABX3 U10410 ( .A(n8225), .B(n8226), .C(n8227), .D(n8228), .Z(
        n8106) );
  HS65_LS_NOR3AX2 U10411 ( .A(n8229), .B(n8230), .C(n8231), .Z(n8228) );
  HS65_LS_NAND4ABX3 U10412 ( .A(n8237), .B(n8238), .C(n8239), .D(n8240), .Z(
        n8225) );
  HS65_LS_NOR4ABX2 U10413 ( .A(n8233), .B(n8234), .C(n8235), .D(n8236), .Z(
        n8227) );
  HS65_LS_NOR4ABX2 U10414 ( .A(n7794), .B(n7795), .C(n7796), .D(n7797), .Z(
        n7699) );
  HS65_LS_NAND4ABX3 U10415 ( .A(n7798), .B(n7799), .C(n7800), .D(n7801), .Z(
        n7797) );
  HS65_LS_NAND4ABX3 U10416 ( .A(n7802), .B(n7803), .C(n7804), .D(n7805), .Z(
        n7796) );
  HS65_LS_AOI222X2 U10417 ( .A(n608), .B(n589), .C(n593), .D(n620), .E(n592), 
        .F(n609), .Z(n7794) );
  HS65_LS_NOR4ABX2 U10418 ( .A(n7894), .B(n7895), .C(n7896), .D(n7897), .Z(
        n7737) );
  HS65_LS_NAND4ABX3 U10419 ( .A(n7898), .B(n7899), .C(n7900), .D(n7901), .Z(
        n7897) );
  HS65_LS_NAND4ABX3 U10420 ( .A(n7902), .B(n7903), .C(n7904), .D(n7905), .Z(
        n7896) );
  HS65_LS_AOI222X2 U10421 ( .A(n121), .B(n102), .C(n106), .D(n133), .E(n105), 
        .F(n122), .Z(n7894) );
  HS65_LS_NOR4ABX2 U10422 ( .A(n7468), .B(n7469), .C(n7470), .D(n7471), .Z(
        n6052) );
  HS65_LS_NAND4ABX3 U10423 ( .A(n6536), .B(n6864), .C(n6343), .D(n6927), .Z(
        n7471) );
  HS65_LS_NAND4ABX3 U10424 ( .A(n6951), .B(n6498), .C(n7475), .D(n6938), .Z(
        n7470) );
  HS65_LS_AOI222X2 U10425 ( .A(n76), .B(n69), .C(n57), .D(n87), .E(n70), .F(
        n74), .Z(n7468) );
  HS65_LS_NOR4ABX2 U10426 ( .A(n5935), .B(n5936), .C(n5937), .D(n5938), .Z(
        n4505) );
  HS65_LS_NAND4ABX3 U10427 ( .A(n4997), .B(n5387), .C(n4789), .D(n5450), .Z(
        n5938) );
  HS65_LS_NAND4ABX3 U10428 ( .A(n5474), .B(n4959), .C(n5942), .D(n5461), .Z(
        n5937) );
  HS65_LS_AOI222X2 U10429 ( .A(n474), .B(n467), .C(n455), .D(n485), .E(n468), 
        .F(n472), .Z(n5935) );
  HS65_LS_NOR4ABX2 U10430 ( .A(n7527), .B(n7528), .C(n7529), .D(n7530), .Z(
        n6098) );
  HS65_LS_NAND4ABX3 U10431 ( .A(n6590), .B(n6979), .C(n6382), .D(n7042), .Z(
        n7530) );
  HS65_LS_NAND4ABX3 U10432 ( .A(n7066), .B(n6552), .C(n7534), .D(n7053), .Z(
        n7529) );
  HS65_LS_AOI222X2 U10433 ( .A(n297), .B(n290), .C(n278), .D(n308), .E(n291), 
        .F(n295), .Z(n7527) );
  HS65_LS_NOR4ABX2 U10434 ( .A(n5876), .B(n5877), .C(n5878), .D(n5879), .Z(
        n4459) );
  HS65_LS_NAND4ABX3 U10435 ( .A(n4943), .B(n5272), .C(n4750), .D(n5335), .Z(
        n5879) );
  HS65_LS_NAND4ABX3 U10436 ( .A(n5359), .B(n4905), .C(n5883), .D(n5346), .Z(
        n5878) );
  HS65_LS_AOI222X2 U10437 ( .A(n255), .B(n248), .C(n236), .D(n266), .E(n249), 
        .F(n253), .Z(n5876) );
  HS65_LS_NOR4ABX2 U10438 ( .A(n5772), .B(n5773), .C(n5774), .D(n5775), .Z(
        n5697) );
  HS65_LS_NAND4ABX3 U10439 ( .A(n4869), .B(n5155), .C(n4643), .D(n5219), .Z(
        n5775) );
  HS65_LS_NAND4ABX3 U10440 ( .A(n5244), .B(n4828), .C(n5776), .D(n5230), .Z(
        n5774) );
  HS65_LS_AOI222X2 U10441 ( .A(n710), .B(n677), .C(n689), .D(n707), .E(n676), 
        .F(n712), .Z(n5772) );
  HS65_LS_NOR4ABX2 U10442 ( .A(n7364), .B(n7365), .C(n7366), .D(n7367), .Z(
        n7289) );
  HS65_LS_NAND4ABX3 U10443 ( .A(n6462), .B(n6747), .C(n6236), .D(n6811), .Z(
        n7367) );
  HS65_LS_NAND4ABX3 U10444 ( .A(n6836), .B(n6421), .C(n7368), .D(n6822), .Z(
        n7366) );
  HS65_LS_AOI222X2 U10445 ( .A(n528), .B(n495), .C(n507), .D(n525), .E(n494), 
        .F(n530), .Z(n7364) );
  HS65_LS_NOR3AX2 U10446 ( .A(n6491), .B(n6515), .C(n6330), .Z(n6853) );
  HS65_LS_NOR3AX2 U10447 ( .A(n4898), .B(n4922), .C(n4737), .Z(n5261) );
  HS65_LS_NOR3AX2 U10448 ( .A(n4952), .B(n4976), .C(n4776), .Z(n5376) );
  HS65_LS_NOR3AX2 U10449 ( .A(n6545), .B(n6569), .C(n6369), .Z(n6968) );
  HS65_LS_NOR3AX2 U10450 ( .A(n4821), .B(n4846), .C(n4629), .Z(n5143) );
  HS65_LS_NOR3AX2 U10451 ( .A(n6414), .B(n6439), .C(n6222), .Z(n6735) );
  HS65_LS_NOR3AX2 U10452 ( .A(n6274), .B(n6299), .C(n6145), .Z(n6614) );
  HS65_LS_NOR3AX2 U10453 ( .A(n4681), .B(n4706), .C(n4552), .Z(n5021) );
  HS65_LS_NAND4ABX3 U10454 ( .A(n3112), .B(n3113), .C(n3114), .D(n3115), .Z(
        n2869) );
  HS65_LS_NOR3X1 U10455 ( .A(n3116), .B(n3117), .C(n3118), .Z(n3115) );
  HS65_LS_AOI222X2 U10456 ( .A(n193), .B(n216), .C(n194), .D(n219), .E(n197), 
        .F(n225), .Z(n3114) );
  HS65_LS_NAND3AX3 U10457 ( .A(n3119), .B(n3120), .C(n3121), .Z(n3113) );
  HS65_LS_NOR3X1 U10458 ( .A(n7868), .B(n8105), .C(n8106), .Z(n8099) );
  HS65_LS_NOR3AX2 U10459 ( .A(n6881), .B(n67), .C(n6865), .Z(n7446) );
  HS65_LS_IVX2 U10460 ( .A(n6344), .Z(n67) );
  HS65_LS_NOR3AX2 U10461 ( .A(n5404), .B(n465), .C(n5388), .Z(n5913) );
  HS65_LS_IVX2 U10462 ( .A(n4790), .Z(n465) );
  HS65_LS_NOR3AX2 U10463 ( .A(n6996), .B(n288), .C(n6980), .Z(n7505) );
  HS65_LS_IVX2 U10464 ( .A(n6383), .Z(n288) );
  HS65_LS_NOR3AX2 U10465 ( .A(n5289), .B(n246), .C(n5273), .Z(n5854) );
  HS65_LS_IVX2 U10466 ( .A(n4751), .Z(n246) );
  HS65_LS_NOR3AX2 U10467 ( .A(n5172), .B(n678), .C(n5156), .Z(n5695) );
  HS65_LS_IVX2 U10468 ( .A(n4644), .Z(n678) );
  HS65_LS_NOR3AX2 U10469 ( .A(n6764), .B(n496), .C(n6748), .Z(n7287) );
  HS65_LS_IVX2 U10470 ( .A(n6237), .Z(n496) );
  HS65_LS_NAND2X2 U10471 ( .A(n395), .B(n365), .Z(n8224) );
  HS65_LS_CBI4I6X2 U10472 ( .A(n81), .B(n83), .C(n61), .D(n6932), .Z(n7209) );
  HS65_LS_CBI4I6X2 U10473 ( .A(n511), .B(n518), .C(n503), .D(n6816), .Z(n7182)
         );
  HS65_LS_CBI4I6X2 U10474 ( .A(n693), .B(n700), .C(n685), .D(n5224), .Z(n5590)
         );
  HS65_LS_CBI4I6X2 U10475 ( .A(n479), .B(n481), .C(n459), .D(n5455), .Z(n5644)
         );
  HS65_LS_CBI4I6X2 U10476 ( .A(n302), .B(n304), .C(n282), .D(n7047), .Z(n7236)
         );
  HS65_LS_CBI4I6X2 U10477 ( .A(n260), .B(n262), .C(n240), .D(n5340), .Z(n5617)
         );
  HS65_LS_NAND4ABX3 U10478 ( .A(n3401), .B(n3402), .C(n3403), .D(n3404), .Z(
        n2999) );
  HS65_LS_NOR3X1 U10479 ( .A(n3405), .B(n3406), .C(n3407), .Z(n3404) );
  HS65_LS_AOI222X2 U10480 ( .A(n419), .B(n441), .C(n422), .D(n443), .E(n420), 
        .F(n434), .Z(n3403) );
  HS65_LS_NAND3AX3 U10481 ( .A(n3408), .B(n3409), .C(n3410), .Z(n3402) );
  HS65_LS_NAND4ABX3 U10482 ( .A(n4307), .B(n4308), .C(n4309), .D(n4310), .Z(
        n3973) );
  HS65_LS_NAND4ABX3 U10483 ( .A(n3408), .B(n3374), .C(n3199), .D(n3387), .Z(
        n4308) );
  HS65_LS_AOI222X2 U10484 ( .A(n438), .B(n424), .C(n440), .D(n415), .E(n437), 
        .F(n413), .Z(n4309) );
  HS65_LS_NAND4ABX3 U10485 ( .A(n3897), .B(n3814), .C(n4311), .D(n3801), .Z(
        n4307) );
  HS65_LS_NAND4ABX3 U10486 ( .A(n4248), .B(n4249), .C(n4250), .D(n4251), .Z(
        n3952) );
  HS65_LS_AOI222X2 U10487 ( .A(n662), .B(n648), .C(n664), .D(n639), .E(n661), 
        .F(n636), .Z(n4250) );
  HS65_LS_NAND4ABX3 U10488 ( .A(n3346), .B(n3312), .C(n3158), .D(n3325), .Z(
        n4249) );
  HS65_LS_NAND4ABX3 U10489 ( .A(n3780), .B(n3697), .C(n4252), .D(n3684), .Z(
        n4248) );
  HS65_LS_NOR2X2 U10490 ( .A(n917), .B(n922), .Z(n2335) );
  HS65_LS_NOR2X2 U10491 ( .A(n835), .B(n840), .Z(n1583) );
  HS65_LS_NOR4ABX2 U10492 ( .A(n6659), .B(n6660), .C(n6661), .D(n6662), .Z(
        n6274) );
  HS65_LS_MX41X4 U10493 ( .D0(n536), .S0(n558), .D1(n568), .S1(n538), .D2(n569), .S2(n542), .D3(n555), .S3(n540), .Z(n6662) );
  HS65_LS_NAND3AX3 U10494 ( .A(n6663), .B(n6664), .C(n6665), .Z(n6661) );
  HS65_LS_NOR4ABX2 U10495 ( .A(n6671), .B(n6672), .C(n6673), .D(n6674), .Z(
        n6659) );
  HS65_LS_NOR4ABX2 U10496 ( .A(n5066), .B(n5067), .C(n5068), .D(n5069), .Z(
        n4681) );
  HS65_LS_MX41X4 U10497 ( .D0(n10), .S0(n32), .D1(n42), .S1(n12), .D2(n43), 
        .S2(n16), .D3(n29), .S3(n14), .Z(n5069) );
  HS65_LS_NAND3AX3 U10498 ( .A(n5070), .B(n5071), .C(n5072), .Z(n5068) );
  HS65_LS_NOR4ABX2 U10499 ( .A(n5078), .B(n5079), .C(n5080), .D(n5081), .Z(
        n5066) );
  HS65_LS_NOR4ABX2 U10500 ( .A(n6896), .B(n6897), .C(n6898), .D(n6899), .Z(
        n6491) );
  HS65_LS_MX41X4 U10501 ( .D0(n68), .S0(n79), .D1(n69), .S1(n91), .D2(n87), 
        .S2(n64), .D3(n81), .S3(n63), .Z(n6899) );
  HS65_LS_NAND3AX3 U10502 ( .A(n6900), .B(n6901), .C(n6902), .Z(n6898) );
  HS65_LS_NOR4ABX2 U10503 ( .A(n6904), .B(n6905), .C(n6906), .D(n6907), .Z(
        n6897) );
  HS65_LS_NOR4ABX2 U10504 ( .A(n5304), .B(n5305), .C(n5306), .D(n5307), .Z(
        n4898) );
  HS65_LS_MX41X4 U10505 ( .D0(n247), .S0(n258), .D1(n248), .S1(n270), .D2(n266), .S2(n243), .D3(n260), .S3(n242), .Z(n5307) );
  HS65_LS_NAND3AX3 U10506 ( .A(n5308), .B(n5309), .C(n5310), .Z(n5306) );
  HS65_LS_NOR4ABX2 U10507 ( .A(n5312), .B(n5313), .C(n5314), .D(n5315), .Z(
        n5305) );
  HS65_LS_NOR4ABX2 U10508 ( .A(n5419), .B(n5420), .C(n5421), .D(n5422), .Z(
        n4952) );
  HS65_LS_MX41X4 U10509 ( .D0(n466), .S0(n477), .D1(n467), .S1(n489), .D2(n485), .S2(n462), .D3(n479), .S3(n461), .Z(n5422) );
  HS65_LS_NAND3AX3 U10510 ( .A(n5423), .B(n5424), .C(n5425), .Z(n5421) );
  HS65_LS_NOR4ABX2 U10511 ( .A(n5427), .B(n5428), .C(n5429), .D(n5430), .Z(
        n5420) );
  HS65_LS_NOR4ABX2 U10512 ( .A(n7011), .B(n7012), .C(n7013), .D(n7014), .Z(
        n6545) );
  HS65_LS_MX41X4 U10513 ( .D0(n289), .S0(n300), .D1(n290), .S1(n312), .D2(n308), .S2(n285), .D3(n302), .S3(n284), .Z(n7014) );
  HS65_LS_NAND3AX3 U10514 ( .A(n7015), .B(n7016), .C(n7017), .Z(n7013) );
  HS65_LS_NOR4ABX2 U10515 ( .A(n7019), .B(n7020), .C(n7021), .D(n7022), .Z(
        n7012) );
  HS65_LS_NOR4ABX2 U10516 ( .A(n5188), .B(n5189), .C(n5190), .D(n5191), .Z(
        n4821) );
  HS65_LS_MX41X4 U10517 ( .D0(n675), .S0(n696), .D1(n677), .S1(n706), .D2(n707), .S2(n681), .D3(n693), .S3(n679), .Z(n5191) );
  HS65_LS_NAND3AX3 U10518 ( .A(n5192), .B(n5193), .C(n5194), .Z(n5190) );
  HS65_LS_NOR4ABX2 U10519 ( .A(n5196), .B(n5197), .C(n5198), .D(n5199), .Z(
        n5189) );
  HS65_LS_NOR4ABX2 U10520 ( .A(n6780), .B(n6781), .C(n6782), .D(n6783), .Z(
        n6414) );
  HS65_LS_MX41X4 U10521 ( .D0(n493), .S0(n514), .D1(n495), .S1(n524), .D2(n525), .S2(n499), .D3(n511), .S3(n497), .Z(n6783) );
  HS65_LS_NAND3AX3 U10522 ( .A(n6784), .B(n6785), .C(n6786), .Z(n6782) );
  HS65_LS_NOR4ABX2 U10523 ( .A(n6788), .B(n6789), .C(n6790), .D(n6791), .Z(
        n6781) );
  HS65_LS_NOR4ABX2 U10524 ( .A(n2464), .B(n2465), .C(n2466), .D(n2467), .Z(
        n2347) );
  HS65_LS_MX41X4 U10525 ( .D0(n923), .S0(n904), .D1(n906), .S1(n917), .D2(n897), .S2(n924), .D3(n895), .S3(n920), .Z(n2467) );
  HS65_LS_NAND3AX3 U10526 ( .A(n2468), .B(n2469), .C(n2470), .Z(n2466) );
  HS65_LS_NOR4ABX2 U10527 ( .A(n2472), .B(n2473), .C(n2474), .D(n2475), .Z(
        n2465) );
  HS65_LS_NOR4ABX2 U10528 ( .A(n1712), .B(n1713), .C(n1714), .D(n1715), .Z(
        n1595) );
  HS65_LS_MX41X4 U10529 ( .D0(n841), .S0(n822), .D1(n824), .S1(n835), .D2(n815), .S2(n842), .D3(n813), .S3(n838), .Z(n1715) );
  HS65_LS_NAND3AX3 U10530 ( .A(n1716), .B(n1717), .C(n1718), .Z(n1714) );
  HS65_LS_NOR4ABX2 U10531 ( .A(n1720), .B(n1721), .C(n1722), .D(n1723), .Z(
        n1713) );
  HS65_LS_NOR4ABX2 U10532 ( .A(n1336), .B(n1337), .C(n1338), .D(n1339), .Z(
        n1219) );
  HS65_LS_MX41X4 U10533 ( .D0(n882), .S0(n863), .D1(n865), .S1(n876), .D2(n856), .S2(n883), .D3(n854), .S3(n879), .Z(n1339) );
  HS65_LS_NAND3AX3 U10534 ( .A(n1340), .B(n1341), .C(n1342), .Z(n1338) );
  HS65_LS_NOR4ABX2 U10535 ( .A(n1344), .B(n1345), .C(n1346), .D(n1347), .Z(
        n1337) );
  HS65_LS_NOR4ABX2 U10536 ( .A(n2088), .B(n2089), .C(n2090), .D(n2091), .Z(
        n1971) );
  HS65_LS_MX41X4 U10537 ( .D0(n800), .S0(n781), .D1(n783), .S1(n794), .D2(n774), .S2(n801), .D3(n772), .S3(n797), .Z(n2091) );
  HS65_LS_NAND3AX3 U10538 ( .A(n2092), .B(n2093), .C(n2094), .Z(n2090) );
  HS65_LS_NOR4ABX2 U10539 ( .A(n2096), .B(n2097), .C(n2098), .D(n2099), .Z(
        n2089) );
  HS65_LS_NOR4ABX2 U10540 ( .A(n3869), .B(n3870), .C(n3871), .D(n3872), .Z(
        n3366) );
  HS65_LS_MX41X4 U10541 ( .D0(n424), .S0(n435), .D1(n445), .S1(n425), .D2(n447), .S2(n420), .D3(n438), .S3(n419), .Z(n3872) );
  HS65_LS_NAND3AX3 U10542 ( .A(n3873), .B(n3874), .C(n3875), .Z(n3871) );
  HS65_LS_NOR4ABX2 U10543 ( .A(n3877), .B(n3878), .C(n3879), .D(n3880), .Z(
        n3870) );
  HS65_LS_NOR4ABX2 U10544 ( .A(n3650), .B(n3651), .C(n3652), .D(n3653), .Z(
        n3237) );
  HS65_LS_NAND4ABX3 U10545 ( .A(n3654), .B(n3655), .C(n3656), .D(n3657), .Z(
        n3652) );
  HS65_LS_MX41X4 U10546 ( .D0(n143), .S0(n167), .D1(n145), .S1(n176), .D2(n177), .S2(n152), .D3(n148), .S3(n165), .Z(n3653) );
  HS65_LS_NOR4ABX2 U10547 ( .A(n3662), .B(n3663), .C(n3664), .D(n3665), .Z(
        n3650) );
  HS65_LS_NOR2X2 U10548 ( .A(n876), .B(n881), .Z(n1207) );
  HS65_LS_NOR2X2 U10549 ( .A(n794), .B(n799), .Z(n1959) );
  HS65_LS_NOR4ABX2 U10550 ( .A(n8717), .B(n8718), .C(n8719), .D(n8720), .Z(
        n8390) );
  HS65_LS_MX41X4 U10551 ( .D0(n591), .S0(n625), .D1(n589), .S1(n618), .D2(n620), .S2(n583), .D3(n623), .S3(n585), .Z(n8720) );
  HS65_LS_NAND3X2 U10552 ( .A(n8721), .B(n7821), .C(n8722), .Z(n8719) );
  HS65_LS_NOR4ABX2 U10553 ( .A(n8724), .B(n7806), .C(n7703), .D(n8725), .Z(
        n8718) );
  HS65_LS_NOR4ABX2 U10554 ( .A(n8805), .B(n8806), .C(n8807), .D(n8808), .Z(
        n8450) );
  HS65_LS_MX41X4 U10555 ( .D0(n104), .S0(n138), .D1(n102), .S1(n131), .D2(n133), .S2(n96), .D3(n136), .S3(n98), .Z(n8808) );
  HS65_LS_NAND3X2 U10556 ( .A(n8809), .B(n7920), .C(n8810), .Z(n8807) );
  HS65_LS_NOR4ABX2 U10557 ( .A(n8812), .B(n7906), .C(n7741), .D(n8813), .Z(
        n8806) );
  HS65_LS_NOR4ABX2 U10558 ( .A(n3752), .B(n3753), .C(n3754), .D(n3755), .Z(
        n3304) );
  HS65_LS_MX41X4 U10559 ( .D0(n648), .S0(n659), .D1(n669), .S1(n649), .D2(n671), .S2(n644), .D3(n662), .S3(n643), .Z(n3755) );
  HS65_LS_NAND3X2 U10560 ( .A(n3756), .B(n3757), .C(n3758), .Z(n3754) );
  HS65_LS_NOR4ABX2 U10561 ( .A(n3760), .B(n3761), .C(n3762), .D(n3763), .Z(
        n3753) );
  HS65_LS_NOR4ABX2 U10562 ( .A(n8290), .B(n8291), .C(n8292), .D(n8293), .Z(
        n8081) );
  HS65_LS_MX41X4 U10563 ( .D0(n402), .S0(n369), .D1(n391), .S1(n367), .D2(n395), .S2(n371), .D3(n370), .S3(n403), .Z(n8293) );
  HS65_LS_NAND3X2 U10564 ( .A(n8294), .B(n8295), .C(n8296), .Z(n8292) );
  HS65_LS_NOR4ABX2 U10565 ( .A(n8302), .B(n8303), .C(n8304), .D(n8305), .Z(
        n8290) );
  HS65_LS_NOR4ABX2 U10566 ( .A(n3511), .B(n3512), .C(n3513), .D(n3514), .Z(
        n3075) );
  HS65_LS_NAND3X2 U10567 ( .A(n3515), .B(n3516), .C(n3517), .Z(n3513) );
  HS65_LS_MX41X4 U10568 ( .D0(n189), .S0(n213), .D1(n223), .S1(n191), .D2(n222), .S2(n197), .D3(n210), .S3(n193), .Z(n3514) );
  HS65_LS_NOR4ABX2 U10569 ( .A(n3519), .B(n3520), .C(n3521), .D(n3522), .Z(
        n3512) );
  HS65_LS_IVX2 U10570 ( .A(n2848), .Z(n415) );
  HS65_LS_IVX2 U10571 ( .A(n2928), .Z(n154) );
  HS65_LS_NOR4ABX2 U10572 ( .A(n8594), .B(n8595), .C(n8596), .D(n8597), .Z(
        n8336) );
  HS65_LS_NAND3AX3 U10573 ( .A(n8598), .B(n8599), .C(n8600), .Z(n8596) );
  HS65_LS_MX41X4 U10574 ( .D0(n343), .S0(n322), .D1(n354), .S1(n319), .D2(n358), .S2(n337), .D3(n335), .S3(n341), .Z(n8597) );
  HS65_LS_NOR4ABX2 U10575 ( .A(n8602), .B(n8603), .C(n8604), .D(n8605), .Z(
        n8595) );
  HS65_LS_NOR3AX2 U10576 ( .A(n1180), .B(n1314), .C(n1351), .Z(n1459) );
  HS65_LS_NOR3AX2 U10577 ( .A(n1932), .B(n2066), .C(n2103), .Z(n2211) );
  HS65_LS_NOR3AX2 U10578 ( .A(n1556), .B(n1690), .C(n1727), .Z(n1835) );
  HS65_LS_NOR3AX2 U10579 ( .A(n2308), .B(n2442), .C(n2479), .Z(n2587) );
  HS65_LS_NOR2X2 U10580 ( .A(n649), .B(n636), .Z(n3352) );
  HS65_LS_IVX2 U10581 ( .A(n7880), .Z(n107) );
  HS65_LS_IVX2 U10582 ( .A(n7817), .Z(n594) );
  HS65_LS_NOR2X2 U10583 ( .A(n425), .B(n413), .Z(n3414) );
  HS65_LS_NOR3AX2 U10584 ( .A(n3196), .B(n3847), .C(n3884), .Z(n4322) );
  HS65_LS_NAND4ABX3 U10585 ( .A(n4139), .B(n4140), .C(n4141), .D(n4142), .Z(
        n3997) );
  HS65_LS_NOR4ABX2 U10586 ( .A(n3582), .B(n3273), .C(n3563), .D(n3598), .Z(
        n4141) );
  HS65_LS_NAND4ABX3 U10587 ( .A(n3269), .B(n3285), .C(n3061), .D(n3048), .Z(
        n4140) );
  HS65_LS_NOR4ABX2 U10588 ( .A(n3629), .B(n3611), .C(n3665), .D(n3637), .Z(
        n4142) );
  HS65_LS_NOR2X2 U10589 ( .A(n77), .B(n84), .Z(n6352) );
  HS65_LS_NOR2X2 U10590 ( .A(n475), .B(n482), .Z(n4798) );
  HS65_LS_NOR2X2 U10591 ( .A(n298), .B(n305), .Z(n6391) );
  HS65_LS_NOR2X2 U10592 ( .A(n256), .B(n263), .Z(n4759) );
  HS65_LS_NOR2X2 U10593 ( .A(n709), .B(n702), .Z(n4652) );
  HS65_LS_NOR2X2 U10594 ( .A(n527), .B(n520), .Z(n6245) );
  HS65_LS_NOR2X2 U10595 ( .A(n45), .B(n38), .Z(n4575) );
  HS65_LS_NOR2X2 U10596 ( .A(n571), .B(n564), .Z(n6168) );
  HS65_LS_NOR2X2 U10597 ( .A(n606), .B(n613), .Z(n7640) );
  HS65_LS_NOR2X2 U10598 ( .A(n119), .B(n126), .Z(n7668) );
  HS65_LS_NOR3X1 U10599 ( .A(n1229), .B(n1230), .C(n1151), .Z(n1222) );
  HS65_LS_NOR3X1 U10600 ( .A(n2357), .B(n2358), .C(n2279), .Z(n2350) );
  HS65_LS_NOR3X1 U10601 ( .A(n1981), .B(n1982), .C(n1903), .Z(n1974) );
  HS65_LS_NOR3X1 U10602 ( .A(n1605), .B(n1606), .C(n1527), .Z(n1598) );
  HS65_LS_NOR2X2 U10603 ( .A(n905), .B(n907), .Z(n2322) );
  HS65_LS_NOR2X2 U10604 ( .A(n823), .B(n825), .Z(n1570) );
  HS65_LS_NOR2X2 U10605 ( .A(n388), .B(n398), .Z(n7997) );
  HS65_LS_NOR2X2 U10606 ( .A(n348), .B(n351), .Z(n8039) );
  HS65_LS_NOR2X2 U10607 ( .A(n864), .B(n866), .Z(n1194) );
  HS65_LS_NOR2X2 U10608 ( .A(n782), .B(n784), .Z(n1946) );
  HS65_LS_NOR2X2 U10609 ( .A(n434), .B(n440), .Z(n3202) );
  HS65_LS_NOR2X2 U10610 ( .A(n225), .B(n217), .Z(n2959) );
  HS65_LS_NOR2X2 U10611 ( .A(n658), .B(n664), .Z(n3161) );
  HS65_LS_NAND4ABX3 U10612 ( .A(n4202), .B(n4203), .C(n4204), .D(n4205), .Z(
        n3935) );
  HS65_LS_NAND4ABX3 U10613 ( .A(n3456), .B(n2968), .C(n3519), .D(n3477), .Z(
        n4203) );
  HS65_LS_NOR4ABX2 U10614 ( .A(n3111), .B(n3496), .C(n3438), .D(n3118), .Z(
        n4205) );
  HS65_LS_MX41X4 U10615 ( .D0(n190), .S0(n213), .D1(n200), .S1(n212), .D2(n219), .S2(n201), .D3(n210), .S3(n198), .Z(n4202) );
  HS65_LS_NOR2X2 U10616 ( .A(n69), .B(n62), .Z(n6480) );
  HS65_LS_NOR2X2 U10617 ( .A(n290), .B(n283), .Z(n6594) );
  HS65_LS_NOR2X2 U10618 ( .A(n248), .B(n241), .Z(n4887) );
  HS65_LS_NOR2X2 U10619 ( .A(n467), .B(n460), .Z(n5001) );
  HS65_LS_NAND4ABX3 U10620 ( .A(n1796), .B(n1797), .C(n1798), .D(n1799), .Z(
        n1773) );
  HS65_LS_NOR4ABX2 U10621 ( .A(n1627), .B(n1698), .C(n1658), .D(n1635), .Z(
        n1799) );
  HS65_LS_NAND4ABX3 U10622 ( .A(n1738), .B(n1565), .C(n1720), .D(n1679), .Z(
        n1797) );
  HS65_LS_NOR4ABX2 U10623 ( .A(n1750), .B(n1730), .C(n1557), .D(n1613), .Z(
        n1798) );
  HS65_LS_NAND4ABX3 U10624 ( .A(n2548), .B(n2549), .C(n2550), .D(n2551), .Z(
        n2525) );
  HS65_LS_NAND4ABX3 U10625 ( .A(n2490), .B(n2317), .C(n2472), .D(n2431), .Z(
        n2549) );
  HS65_LS_NOR4ABX2 U10626 ( .A(n2379), .B(n2450), .C(n2410), .D(n2387), .Z(
        n2551) );
  HS65_LS_NOR4ABX2 U10627 ( .A(n2502), .B(n2482), .C(n2309), .D(n2365), .Z(
        n2550) );
  HS65_LS_NAND4ABX3 U10628 ( .A(n1420), .B(n1421), .C(n1422), .D(n1423), .Z(
        n1397) );
  HS65_LS_NAND4ABX3 U10629 ( .A(n1362), .B(n1189), .C(n1344), .D(n1303), .Z(
        n1421) );
  HS65_LS_NOR4ABX2 U10630 ( .A(n1251), .B(n1322), .C(n1282), .D(n1259), .Z(
        n1423) );
  HS65_LS_NOR4ABX2 U10631 ( .A(n1374), .B(n1354), .C(n1181), .D(n1237), .Z(
        n1422) );
  HS65_LS_NAND4ABX3 U10632 ( .A(n2172), .B(n2173), .C(n2174), .D(n2175), .Z(
        n2149) );
  HS65_LS_NAND4ABX3 U10633 ( .A(n2114), .B(n1941), .C(n2096), .D(n2055), .Z(
        n2173) );
  HS65_LS_NOR4ABX2 U10634 ( .A(n2003), .B(n2074), .C(n2034), .D(n2011), .Z(
        n2175) );
  HS65_LS_NOR4ABX2 U10635 ( .A(n2126), .B(n2106), .C(n1933), .D(n1989), .Z(
        n2174) );
  HS65_LS_NOR3X1 U10636 ( .A(n7971), .B(n8401), .C(n8402), .Z(n8394) );
  HS65_LS_NOR3X1 U10637 ( .A(n7984), .B(n8461), .C(n8462), .Z(n8454) );
  HS65_LS_NOR3X1 U10638 ( .A(n3248), .B(n3249), .C(n2920), .Z(n3241) );
  HS65_LS_NOR3X1 U10639 ( .A(n3086), .B(n3087), .C(n2870), .Z(n3079) );
  HS65_LS_NOR3X1 U10640 ( .A(n3377), .B(n3378), .C(n3000), .Z(n3370) );
  HS65_LS_NOR3X1 U10641 ( .A(n3315), .B(n3316), .C(n2982), .Z(n3308) );
  HS65_LS_NOR3X1 U10642 ( .A(n3619), .B(n3037), .C(n3654), .Z(n4106) );
  HS65_LS_NAND2X2 U10643 ( .A(n403), .B(n365), .Z(n8270) );
  HS65_LS_NOR4ABX2 U10644 ( .A(n4076), .B(n4077), .C(n4078), .D(n4079), .Z(
        n3906) );
  HS65_LS_NAND4ABX3 U10645 ( .A(n3430), .B(n3084), .C(n4080), .D(n3443), .Z(
        n4079) );
  HS65_LS_MX41X4 U10646 ( .D0(n190), .S0(n210), .D1(n222), .S1(n201), .D2(n223), .S2(n198), .D3(n199), .S3(n215), .Z(n4078) );
  HS65_LS_AOI222X2 U10647 ( .A(n221), .B(n191), .C(n200), .D(n226), .E(n219), 
        .F(n205), .Z(n4076) );
  HS65_LS_NAND4ABX3 U10648 ( .A(n3031), .B(n3032), .C(n3033), .D(n3034), .Z(
        n2919) );
  HS65_LS_NOR3AX2 U10649 ( .A(n3039), .B(n3040), .C(n3041), .Z(n3033) );
  HS65_LS_NOR4ABX2 U10650 ( .A(n3035), .B(n3036), .C(n3037), .D(n3038), .Z(
        n3034) );
  HS65_LS_NAND3AX3 U10651 ( .A(n3047), .B(n3048), .C(n3049), .Z(n3031) );
  HS65_LS_NOR4ABX2 U10652 ( .A(n9045), .B(n9046), .C(n9047), .D(n9048), .Z(
        n7688) );
  HS65_LS_NAND4ABX3 U10653 ( .A(n8682), .B(n8702), .C(n8397), .D(n9049), .Z(
        n9048) );
  HS65_LS_MX41X4 U10654 ( .D0(n623), .S0(n592), .D1(n596), .S1(n620), .D2(n597), .S2(n618), .D3(n612), .S3(n594), .Z(n9047) );
  HS65_LS_NOR4ABX2 U10655 ( .A(n8726), .B(n8716), .C(n8410), .D(n8763), .Z(
        n9046) );
  HS65_LS_NOR4ABX2 U10656 ( .A(n9103), .B(n9104), .C(n9105), .D(n9106), .Z(
        n7726) );
  HS65_LS_NAND4ABX3 U10657 ( .A(n8770), .B(n8790), .C(n8457), .D(n9107), .Z(
        n9106) );
  HS65_LS_MX41X4 U10658 ( .D0(n136), .S0(n105), .D1(n109), .S1(n133), .D2(n110), .S2(n131), .D3(n125), .S3(n107), .Z(n9105) );
  HS65_LS_NOR4ABX2 U10659 ( .A(n8814), .B(n8804), .C(n8470), .D(n8851), .Z(
        n9104) );
  HS65_LS_NOR4ABX2 U10660 ( .A(n8659), .B(n8660), .C(n8661), .D(n8662), .Z(
        n7763) );
  HS65_LS_NAND4ABX3 U10661 ( .A(n8089), .B(n8245), .C(n8312), .D(n8111), .Z(
        n8662) );
  HS65_LS_NAND4ABX3 U10662 ( .A(n8261), .B(n8022), .C(n8223), .D(n8276), .Z(
        n8661) );
  HS65_LS_NOR4ABX2 U10663 ( .A(n8664), .B(n8128), .C(n8301), .D(n8235), .Z(
        n8660) );
  HS65_LS_NOR4ABX2 U10664 ( .A(n8868), .B(n8869), .C(n8870), .D(n8871), .Z(
        n7780) );
  HS65_LS_NAND4ABX3 U10665 ( .A(n8383), .B(n8549), .C(n8539), .D(n8353), .Z(
        n8871) );
  HS65_LS_NOR4ABX2 U10666 ( .A(n8872), .B(n8370), .C(n8605), .D(n8614), .Z(
        n8869) );
  HS65_LS_NAND4ABX3 U10667 ( .A(n8565), .B(n8527), .C(n8065), .D(n8580), .Z(
        n8870) );
  HS65_LS_NOR4ABX2 U10668 ( .A(n9025), .B(n9026), .C(n9027), .D(n9028), .Z(
        n7636) );
  HS65_LS_NAND4ABX3 U10669 ( .A(n8166), .B(n8738), .C(n8727), .D(n8697), .Z(
        n9028) );
  HS65_LS_NOR4ABX2 U10670 ( .A(n8746), .B(n8411), .C(n8730), .D(n8158), .Z(
        n9025) );
  HS65_LS_MX41X4 U10671 ( .D0(n592), .S0(n625), .D1(n593), .S1(n624), .D2(n596), .S2(n616), .D3(n623), .S3(n597), .Z(n9027) );
  HS65_LS_NOR4ABX2 U10672 ( .A(n9083), .B(n9084), .C(n9085), .D(n9086), .Z(
        n7664) );
  HS65_LS_NAND4ABX3 U10673 ( .A(n8198), .B(n8826), .C(n8815), .D(n8785), .Z(
        n9086) );
  HS65_LS_NOR4ABX2 U10674 ( .A(n8834), .B(n8471), .C(n8818), .D(n8190), .Z(
        n9083) );
  HS65_LS_MX41X4 U10675 ( .D0(n105), .S0(n138), .D1(n106), .S1(n137), .D2(n109), .S2(n129), .D3(n136), .S3(n110), .Z(n9085) );
  HS65_LS_CBI4I6X2 U10676 ( .A(n165), .B(n171), .C(n160), .D(n3577), .Z(n4003)
         );
  HS65_LS_NOR4ABX2 U10677 ( .A(n3600), .B(n3601), .C(n3602), .D(n3603), .Z(
        n2917) );
  HS65_LS_NAND4ABX3 U10678 ( .A(n3604), .B(n3605), .C(n3606), .D(n3607), .Z(
        n3603) );
  HS65_LS_MX41X4 U10679 ( .D0(n149), .S0(n167), .D1(n155), .S1(n174), .D2(n145), .S2(n166), .D3(n160), .S3(n3608), .Z(n3602) );
  HS65_LS_AOI212X2 U10680 ( .A(n168), .B(n3609), .C(n152), .D(n3234), .E(n3610), .Z(n3601) );
  HS65_LS_NOR4ABX2 U10681 ( .A(n5904), .B(n5905), .C(n5906), .D(n5907), .Z(
        n5561) );
  HS65_LS_NAND4ABX3 U10682 ( .A(n5435), .B(n4988), .C(n4962), .D(n5456), .Z(
        n5907) );
  HS65_LS_NAND4ABX3 U10683 ( .A(n4795), .B(n5411), .C(n5398), .D(n5449), .Z(
        n5906) );
  HS65_LS_AOI222X2 U10684 ( .A(n467), .B(n481), .C(n459), .D(n478), .E(n489), 
        .F(n457), .Z(n5904) );
  HS65_LS_NOR4ABX2 U10685 ( .A(n5845), .B(n5846), .C(n5847), .D(n5848), .Z(
        n5540) );
  HS65_LS_NAND4ABX3 U10686 ( .A(n5320), .B(n4934), .C(n4908), .D(n5341), .Z(
        n5848) );
  HS65_LS_NAND4ABX3 U10687 ( .A(n4756), .B(n5296), .C(n5283), .D(n5334), .Z(
        n5847) );
  HS65_LS_AOI222X2 U10688 ( .A(n248), .B(n262), .C(n240), .D(n259), .E(n270), 
        .F(n238), .Z(n5845) );
  HS65_LS_NOR4ABX2 U10689 ( .A(n7496), .B(n7497), .C(n7498), .D(n7499), .Z(
        n7153) );
  HS65_LS_NAND4ABX3 U10690 ( .A(n7027), .B(n6581), .C(n6555), .D(n7048), .Z(
        n7499) );
  HS65_LS_NAND4ABX3 U10691 ( .A(n6388), .B(n7003), .C(n6990), .D(n7041), .Z(
        n7498) );
  HS65_LS_AOI222X2 U10692 ( .A(n290), .B(n304), .C(n282), .D(n301), .E(n312), 
        .F(n280), .Z(n7496) );
  HS65_LS_NOR4ABX2 U10693 ( .A(n5805), .B(n5806), .C(n5807), .D(n5808), .Z(
        n5684) );
  HS65_LS_NAND4ABX3 U10694 ( .A(n5204), .B(n4858), .C(n4831), .D(n5225), .Z(
        n5808) );
  HS65_LS_NAND4ABX3 U10695 ( .A(n4649), .B(n5179), .C(n5166), .D(n5218), .Z(
        n5807) );
  HS65_LS_AOI222X2 U10696 ( .A(n677), .B(n700), .C(n685), .D(n697), .E(n706), 
        .F(n684), .Z(n5805) );
  HS65_LS_NOR4ABX2 U10697 ( .A(n5743), .B(n5744), .C(n5745), .D(n5746), .Z(
        n5654) );
  HS65_LS_NAND4ABX3 U10698 ( .A(n5082), .B(n4718), .C(n4691), .D(n5119), .Z(
        n5746) );
  HS65_LS_NAND4ABX3 U10699 ( .A(n5057), .B(n4572), .C(n5044), .D(n5096), .Z(
        n5745) );
  HS65_LS_AOI222X2 U10700 ( .A(n12), .B(n36), .C(n21), .D(n33), .E(n42), .F(
        n20), .Z(n5743) );
  HS65_LS_NOR4ABX2 U10701 ( .A(n7397), .B(n7398), .C(n7399), .D(n7400), .Z(
        n7276) );
  HS65_LS_NAND4ABX3 U10702 ( .A(n6796), .B(n6451), .C(n6424), .D(n6817), .Z(
        n7400) );
  HS65_LS_NAND4ABX3 U10703 ( .A(n6242), .B(n6771), .C(n6758), .D(n6810), .Z(
        n7399) );
  HS65_LS_AOI222X2 U10704 ( .A(n495), .B(n518), .C(n503), .D(n515), .E(n524), 
        .F(n502), .Z(n7397) );
  HS65_LS_NOR4ABX2 U10705 ( .A(n7437), .B(n7438), .C(n7439), .D(n7440), .Z(
        n7132) );
  HS65_LS_NAND4ABX3 U10706 ( .A(n6912), .B(n6527), .C(n6501), .D(n6933), .Z(
        n7440) );
  HS65_LS_NAND4ABX3 U10707 ( .A(n6349), .B(n6888), .C(n6875), .D(n6926), .Z(
        n7439) );
  HS65_LS_AOI222X2 U10708 ( .A(n69), .B(n83), .C(n61), .D(n80), .E(n91), .F(
        n59), .Z(n7437) );
  HS65_LS_NOR4ABX2 U10709 ( .A(n7335), .B(n7336), .C(n7337), .D(n7338), .Z(
        n7246) );
  HS65_LS_NAND4ABX3 U10710 ( .A(n6675), .B(n6311), .C(n6284), .D(n6712), .Z(
        n7338) );
  HS65_LS_NAND4ABX3 U10711 ( .A(n6650), .B(n6165), .C(n6637), .D(n6689), .Z(
        n7337) );
  HS65_LS_AOI222X2 U10712 ( .A(n538), .B(n562), .C(n547), .D(n559), .E(n568), 
        .F(n546), .Z(n7335) );
  HS65_LS_NAND2X2 U10713 ( .A(n61), .B(n76), .Z(n6538) );
  HS65_LS_NAND2X2 U10714 ( .A(n282), .B(n297), .Z(n6592) );
  HS65_LS_NAND2X2 U10715 ( .A(n459), .B(n474), .Z(n4999) );
  HS65_LS_NAND2X2 U10716 ( .A(n240), .B(n255), .Z(n4945) );
  HS65_LS_NAND2X2 U10717 ( .A(n685), .B(n710), .Z(n4871) );
  HS65_LS_NAND2X2 U10718 ( .A(n503), .B(n528), .Z(n6464) );
  HS65_LS_NOR4ABX2 U10719 ( .A(n8990), .B(n8991), .C(n8992), .D(n8993), .Z(
        n8656) );
  HS65_LS_NAND4ABX3 U10720 ( .A(n8222), .B(n8006), .C(n8299), .D(n8259), .Z(
        n8993) );
  HS65_LS_MX41X4 U10721 ( .D0(n366), .S0(n402), .D1(n381), .S1(n404), .D2(n393), .S2(n379), .D3(n403), .S3(n380), .Z(n8992) );
  HS65_LS_NOR4ABX2 U10722 ( .A(n8127), .B(n8087), .C(n8278), .D(n8236), .Z(
        n8991) );
  HS65_LS_NAND4ABX3 U10723 ( .A(n3431), .B(n3432), .C(n3433), .D(n3434), .Z(
        n3086) );
  HS65_LS_NAND3X2 U10724 ( .A(n3443), .B(n3444), .C(n3445), .Z(n3431) );
  HS65_LS_NOR4ABX2 U10725 ( .A(n3439), .B(n3440), .C(n3441), .D(n3442), .Z(
        n3433) );
  HS65_LS_NOR4ABX2 U10726 ( .A(n3435), .B(n3436), .C(n3437), .D(n3438), .Z(
        n3434) );
  HS65_LS_NOR4ABX2 U10727 ( .A(n4019), .B(n4020), .C(n4021), .D(n4022), .Z(
        n3959) );
  HS65_LS_NAND4ABX3 U10728 ( .A(n3720), .B(n3170), .C(n3700), .D(n3760), .Z(
        n4022) );
  HS65_LS_MX41X4 U10729 ( .D0(n650), .S0(n659), .D1(n641), .S1(n661), .D2(n667), .S2(n640), .D3(n662), .S3(n637), .Z(n4021) );
  HS65_LS_NOR4ABX2 U10730 ( .A(n3337), .B(n3738), .C(n3682), .D(n3345), .Z(
        n4020) );
  HS65_LS_NOR4ABX2 U10731 ( .A(n8241), .B(n8242), .C(n8243), .D(n8244), .Z(
        n7873) );
  HS65_LS_NAND4ABX3 U10732 ( .A(n8245), .B(n8246), .C(n8247), .D(n8248), .Z(
        n8244) );
  HS65_LS_MX41X4 U10733 ( .D0(n372), .S0(n402), .D1(n393), .S1(n381), .D2(n404), .S2(n367), .D3(n375), .S3(n8249), .Z(n8243) );
  HS65_LS_AOI212X2 U10734 ( .A(n401), .B(n8250), .C(n371), .D(n8078), .E(n8251), .Z(n8242) );
  HS65_LS_NOR4ABX2 U10735 ( .A(n4043), .B(n4044), .C(n4045), .D(n4046), .Z(
        n3980) );
  HS65_LS_NAND4ABX3 U10736 ( .A(n3816), .B(n3211), .C(n3877), .D(n3836), .Z(
        n4046) );
  HS65_LS_MX41X4 U10737 ( .D0(n426), .S0(n435), .D1(n417), .S1(n437), .D2(n443), .S2(n416), .D3(n438), .S3(n414), .Z(n4045) );
  HS65_LS_NOR4ABX2 U10738 ( .A(n3400), .B(n3855), .C(n3799), .D(n3407), .Z(
        n4044) );
  HS65_LS_NAND2X2 U10739 ( .A(n550), .B(n572), .Z(n6611) );
  HS65_LS_NAND2X2 U10740 ( .A(n24), .B(n46), .Z(n5018) );
  HS65_LS_NAND4ABX3 U10741 ( .A(n3675), .B(n3676), .C(n3677), .D(n3678), .Z(
        n3315) );
  HS65_LS_NAND3X2 U10742 ( .A(n3687), .B(n3688), .C(n3689), .Z(n3675) );
  HS65_LS_NOR4ABX2 U10743 ( .A(n3683), .B(n3684), .C(n3685), .D(n3686), .Z(
        n3677) );
  HS65_LS_NOR4ABX2 U10744 ( .A(n3679), .B(n3680), .C(n3681), .D(n3682), .Z(
        n3678) );
  HS65_LS_NAND2X2 U10745 ( .A(n21), .B(n46), .Z(n4731) );
  HS65_LS_NAND2X2 U10746 ( .A(n547), .B(n572), .Z(n6324) );
  HS65_LS_NAND4ABX3 U10747 ( .A(n2403), .B(n2404), .C(n2405), .D(n2406), .Z(
        n2357) );
  HS65_LS_NAND3X2 U10748 ( .A(n2415), .B(n2416), .C(n2417), .Z(n2403) );
  HS65_LS_NOR4ABX2 U10749 ( .A(n2407), .B(n2408), .C(n2409), .D(n2410), .Z(
        n2406) );
  HS65_LS_NOR4ABX2 U10750 ( .A(n2411), .B(n2412), .C(n2413), .D(n2414), .Z(
        n2405) );
  HS65_LS_NAND4ABX3 U10751 ( .A(n1651), .B(n1652), .C(n1653), .D(n1654), .Z(
        n1605) );
  HS65_LS_NAND3X2 U10752 ( .A(n1663), .B(n1664), .C(n1665), .Z(n1651) );
  HS65_LS_NOR4ABX2 U10753 ( .A(n1655), .B(n1656), .C(n1657), .D(n1658), .Z(
        n1654) );
  HS65_LS_NOR4ABX2 U10754 ( .A(n1659), .B(n1660), .C(n1661), .D(n1662), .Z(
        n1653) );
  HS65_LS_NAND4ABX3 U10755 ( .A(n1275), .B(n1276), .C(n1277), .D(n1278), .Z(
        n1229) );
  HS65_LS_NAND3X2 U10756 ( .A(n1287), .B(n1288), .C(n1289), .Z(n1275) );
  HS65_LS_NOR4ABX2 U10757 ( .A(n1279), .B(n1280), .C(n1281), .D(n1282), .Z(
        n1278) );
  HS65_LS_NOR4ABX2 U10758 ( .A(n1283), .B(n1284), .C(n1285), .D(n1286), .Z(
        n1277) );
  HS65_LS_NAND4ABX3 U10759 ( .A(n3792), .B(n3793), .C(n3794), .D(n3795), .Z(
        n3377) );
  HS65_LS_NOR4ABX2 U10760 ( .A(n3796), .B(n3797), .C(n3798), .D(n3799), .Z(
        n3795) );
  HS65_LS_NOR4ABX2 U10761 ( .A(n3800), .B(n3801), .C(n3802), .D(n3803), .Z(
        n3794) );
  HS65_LS_NAND3X2 U10762 ( .A(n3804), .B(n3805), .C(n3806), .Z(n3792) );
  HS65_LS_NAND4ABX3 U10763 ( .A(n2027), .B(n2028), .C(n2029), .D(n2030), .Z(
        n1981) );
  HS65_LS_NAND3X2 U10764 ( .A(n2039), .B(n2040), .C(n2041), .Z(n2027) );
  HS65_LS_NOR4ABX2 U10765 ( .A(n2031), .B(n2032), .C(n2033), .D(n2034), .Z(
        n2030) );
  HS65_LS_NOR4ABX2 U10766 ( .A(n2035), .B(n2036), .C(n2037), .D(n2038), .Z(
        n2029) );
  HS65_LS_NAND4ABX3 U10767 ( .A(n3557), .B(n3558), .C(n3559), .D(n3560), .Z(
        n3248) );
  HS65_LS_NOR4ABX2 U10768 ( .A(n3565), .B(n3566), .C(n3567), .D(n3568), .Z(
        n3559) );
  HS65_LS_NAND3AX3 U10769 ( .A(n3569), .B(n3570), .C(n3571), .Z(n3557) );
  HS65_LS_NOR4ABX2 U10770 ( .A(n3561), .B(n3562), .C(n3563), .D(n3564), .Z(
        n3560) );
  HS65_LS_NAND2X2 U10771 ( .A(n388), .B(n367), .Z(n8276) );
  HS65_LS_NAND2X2 U10772 ( .A(n348), .B(n319), .Z(n8580) );
  HS65_LS_NOR4ABX2 U10773 ( .A(n5739), .B(n5740), .C(n5741), .D(n5742), .Z(
        n5513) );
  HS65_LS_NAND4ABX3 U10774 ( .A(n5093), .B(n4584), .C(n5071), .D(n5045), .Z(
        n5742) );
  HS65_LS_MX41X4 U10775 ( .D0(n11), .S0(n32), .D1(n25), .S1(n31), .D2(n40), 
        .S2(n26), .D3(n29), .S3(n23), .Z(n5741) );
  HS65_LS_NOR4ABX2 U10776 ( .A(n4690), .B(n5103), .C(n4704), .D(n5062), .Z(
        n5740) );
  HS65_LS_NOR4ABX2 U10777 ( .A(n7331), .B(n7332), .C(n7333), .D(n7334), .Z(
        n7105) );
  HS65_LS_NAND4ABX3 U10778 ( .A(n6686), .B(n6177), .C(n6664), .D(n6638), .Z(
        n7334) );
  HS65_LS_MX41X4 U10779 ( .D0(n537), .S0(n558), .D1(n551), .S1(n557), .D2(n566), .S2(n552), .D3(n555), .S3(n549), .Z(n7333) );
  HS65_LS_NOR4ABX2 U10780 ( .A(n6283), .B(n6696), .C(n6297), .D(n6655), .Z(
        n7332) );
  HS65_LS_NAND2X2 U10781 ( .A(n586), .B(n624), .Z(n8413) );
  HS65_LS_NAND2X2 U10782 ( .A(n99), .B(n137), .Z(n8473) );
  HS65_LS_NOR4ABX2 U10783 ( .A(n5635), .B(n5636), .C(n5637), .D(n5638), .Z(
        n5562) );
  HS65_LS_NAND4ABX3 U10784 ( .A(n4807), .B(n5446), .C(n5399), .D(n5424), .Z(
        n5638) );
  HS65_LS_MX41X4 U10785 ( .D0(n468), .S0(n477), .D1(n455), .S1(n480), .D2(n487), .S2(n456), .D3(n479), .S3(n453), .Z(n5637) );
  HS65_LS_NOR4ABX2 U10786 ( .A(n4961), .B(n5469), .C(n4974), .D(n5415), .Z(
        n5636) );
  HS65_LS_NOR4ABX2 U10787 ( .A(n5608), .B(n5609), .C(n5610), .D(n5611), .Z(
        n5541) );
  HS65_LS_NAND4ABX3 U10788 ( .A(n4768), .B(n5331), .C(n5284), .D(n5309), .Z(
        n5611) );
  HS65_LS_MX41X4 U10789 ( .D0(n249), .S0(n258), .D1(n236), .S1(n261), .D2(n268), .S2(n237), .D3(n260), .S3(n234), .Z(n5610) );
  HS65_LS_NOR4ABX2 U10790 ( .A(n4907), .B(n5354), .C(n4920), .D(n5300), .Z(
        n5609) );
  HS65_LS_NOR4ABX2 U10791 ( .A(n7227), .B(n7228), .C(n7229), .D(n7230), .Z(
        n7154) );
  HS65_LS_NAND4ABX3 U10792 ( .A(n6400), .B(n7038), .C(n6991), .D(n7016), .Z(
        n7230) );
  HS65_LS_MX41X4 U10793 ( .D0(n291), .S0(n300), .D1(n278), .S1(n303), .D2(n310), .S2(n279), .D3(n302), .S3(n276), .Z(n7229) );
  HS65_LS_NOR4ABX2 U10794 ( .A(n6554), .B(n7061), .C(n6567), .D(n7007), .Z(
        n7228) );
  HS65_LS_NOR4ABX2 U10795 ( .A(n5801), .B(n5802), .C(n5803), .D(n5804), .Z(
        n5578) );
  HS65_LS_NAND4ABX3 U10796 ( .A(n4661), .B(n5215), .C(n5167), .D(n5193), .Z(
        n5804) );
  HS65_LS_MX41X4 U10797 ( .D0(n676), .S0(n696), .D1(n689), .S1(n695), .D2(n704), .S2(n690), .D3(n693), .S3(n687), .Z(n5803) );
  HS65_LS_NOR4ABX2 U10798 ( .A(n4830), .B(n5239), .C(n4844), .D(n5184), .Z(
        n5802) );
  HS65_LS_NOR4ABX2 U10799 ( .A(n7393), .B(n7394), .C(n7395), .D(n7396), .Z(
        n7170) );
  HS65_LS_NAND4ABX3 U10800 ( .A(n6254), .B(n6807), .C(n6759), .D(n6785), .Z(
        n7396) );
  HS65_LS_MX41X4 U10801 ( .D0(n494), .S0(n514), .D1(n507), .S1(n513), .D2(n522), .S2(n508), .D3(n511), .S3(n505), .Z(n7395) );
  HS65_LS_NOR4ABX2 U10802 ( .A(n6423), .B(n6831), .C(n6437), .D(n6776), .Z(
        n7394) );
  HS65_LS_NOR4ABX2 U10803 ( .A(n7200), .B(n7201), .C(n7202), .D(n7203), .Z(
        n7133) );
  HS65_LS_NAND4ABX3 U10804 ( .A(n6361), .B(n6923), .C(n6876), .D(n6901), .Z(
        n7203) );
  HS65_LS_MX41X4 U10805 ( .D0(n70), .S0(n79), .D1(n57), .S1(n82), .D2(n89), 
        .S2(n58), .D3(n81), .S3(n55), .Z(n7202) );
  HS65_LS_NOR4ABX2 U10806 ( .A(n6500), .B(n6946), .C(n6513), .D(n6892), .Z(
        n7201) );
  HS65_LS_NOR4ABX2 U10807 ( .A(n9020), .B(n9021), .C(n9022), .D(n9023), .Z(
        n7689) );
  HS65_LS_NAND4ABX3 U10808 ( .A(n8715), .B(n8737), .C(n8703), .D(n8152), .Z(
        n9022) );
  HS65_LS_NAND4ABX3 U10809 ( .A(n8426), .B(n8745), .C(n8690), .D(n8413), .Z(
        n9023) );
  HS65_LS_AOI222X2 U10810 ( .A(n589), .B(n615), .C(n622), .D(n601), .E(n600), 
        .F(n618), .Z(n9020) );
  HS65_LS_NOR4ABX2 U10811 ( .A(n9078), .B(n9079), .C(n9080), .D(n9081), .Z(
        n7727) );
  HS65_LS_NAND4ABX3 U10812 ( .A(n8803), .B(n8825), .C(n8791), .D(n8184), .Z(
        n9080) );
  HS65_LS_NAND4ABX3 U10813 ( .A(n8486), .B(n8833), .C(n8778), .D(n8473), .Z(
        n9081) );
  HS65_LS_AOI222X2 U10814 ( .A(n102), .B(n128), .C(n135), .D(n114), .E(n113), 
        .F(n131), .Z(n9078) );
  HS65_LS_NOR4ABX2 U10815 ( .A(n4328), .B(n4329), .C(n4330), .D(n4331), .Z(
        n3971) );
  HS65_LS_NAND4ABX3 U10816 ( .A(n3791), .B(n3375), .C(n4332), .D(n3804), .Z(
        n4331) );
  HS65_LS_MX41X4 U10817 ( .D0(n426), .S0(n438), .D1(n447), .S1(n416), .D2(n445), .S2(n414), .D3(n415), .S3(n442), .Z(n4330) );
  HS65_LS_AOI222X2 U10818 ( .A(n446), .B(n425), .C(n417), .D(n432), .E(n443), 
        .F(n411), .Z(n4328) );
  HS65_LS_NOR4ABX2 U10819 ( .A(n4269), .B(n4270), .C(n4271), .D(n4272), .Z(
        n3950) );
  HS65_LS_NAND4ABX3 U10820 ( .A(n3674), .B(n3313), .C(n4273), .D(n3687), .Z(
        n4272) );
  HS65_LS_MX41X4 U10821 ( .D0(n650), .S0(n662), .D1(n671), .S1(n640), .D2(n669), .S2(n637), .D3(n639), .S3(n666), .Z(n4271) );
  HS65_LS_AOI222X2 U10822 ( .A(n670), .B(n649), .C(n641), .D(n656), .E(n667), 
        .F(n634), .Z(n4269) );
  HS65_LS_NOR4ABX2 U10823 ( .A(n3819), .B(n3820), .C(n3821), .D(n3822), .Z(
        n2997) );
  HS65_LS_NAND4ABX3 U10824 ( .A(n3823), .B(n3824), .C(n3825), .D(n3826), .Z(
        n3822) );
  HS65_LS_MX41X4 U10825 ( .D0(n422), .S0(n435), .D1(n443), .S1(n417), .D2(n437), .S2(n425), .D3(n411), .S3(n3827), .Z(n3821) );
  HS65_LS_AOI212X2 U10826 ( .A(n436), .B(n3828), .C(n420), .D(n3364), .E(n3829), .Z(n3820) );
  HS65_LS_NOR4ABX2 U10827 ( .A(n3459), .B(n3460), .C(n3461), .D(n3462), .Z(
        n2867) );
  HS65_LS_MX41X4 U10828 ( .D0(n194), .S0(n213), .D1(n219), .S1(n200), .D2(n212), .S2(n191), .D3(n205), .S3(n3467), .Z(n3461) );
  HS65_LS_NAND4ABX3 U10829 ( .A(n3463), .B(n3464), .C(n3465), .D(n3466), .Z(
        n3462) );
  HS65_LS_AOI212X2 U10830 ( .A(n214), .B(n3468), .C(n197), .D(n3072), .E(n3469), .Z(n3460) );
  HS65_LS_NOR4ABX2 U10831 ( .A(n3702), .B(n3703), .C(n3704), .D(n3705), .Z(
        n2979) );
  HS65_LS_NAND4ABX3 U10832 ( .A(n3706), .B(n3707), .C(n3708), .D(n3709), .Z(
        n3705) );
  HS65_LS_MX41X4 U10833 ( .D0(n646), .S0(n659), .D1(n667), .S1(n641), .D2(n661), .S2(n649), .D3(n634), .S3(n3710), .Z(n3704) );
  HS65_LS_AOI212X2 U10834 ( .A(n660), .B(n3711), .C(n644), .D(n3302), .E(n3712), .Z(n3703) );
  HS65_LS_NOR4ABX2 U10835 ( .A(n4143), .B(n4144), .C(n4145), .D(n4146), .Z(
        n4091) );
  HS65_LS_OR4X4 U10836 ( .A(n3640), .B(n3660), .C(n3621), .D(n3604), .Z(n4145)
         );
  HS65_LS_NAND4ABX3 U10837 ( .A(n3288), .B(n3245), .C(n3036), .D(n3259), .Z(
        n4146) );
  HS65_LS_AOI222X2 U10838 ( .A(n145), .B(n171), .C(n160), .D(n168), .E(n158), 
        .F(n176), .Z(n4143) );
  HS65_LS_NOR4ABX2 U10839 ( .A(n8922), .B(n8923), .C(n8924), .D(n8925), .Z(
        n8865) );
  HS65_LS_NAND4ABX3 U10840 ( .A(n8604), .B(n8048), .C(n8528), .D(n8563), .Z(
        n8925) );
  HS65_LS_MX41X4 U10841 ( .D0(n321), .S0(n343), .D1(n332), .S1(n345), .D2(n357), .S2(n330), .D3(n341), .S3(n331), .Z(n8924) );
  HS65_LS_NOR4ABX2 U10842 ( .A(n8540), .B(n8551), .C(n8064), .D(n8355), .Z(
        n8922) );
  HS65_LS_NOR4ABX2 U10843 ( .A(n1846), .B(n1847), .C(n1848), .D(n1849), .Z(
        n1772) );
  HS65_LS_NAND4ABX3 U10844 ( .A(n1558), .B(n1681), .C(n1740), .D(n1697), .Z(
        n1848) );
  HS65_LS_NAND4ABX3 U10845 ( .A(n1634), .B(n1728), .C(n1749), .D(n1611), .Z(
        n1849) );
  HS65_LS_AOI222X2 U10846 ( .A(n821), .B(n835), .C(n817), .D(n847), .E(n833), 
        .F(n824), .Z(n1846) );
  HS65_LS_NOR4ABX2 U10847 ( .A(n2598), .B(n2599), .C(n2600), .D(n2601), .Z(
        n2524) );
  HS65_LS_NAND4ABX3 U10848 ( .A(n2310), .B(n2433), .C(n2492), .D(n2449), .Z(
        n2600) );
  HS65_LS_NAND4ABX3 U10849 ( .A(n2386), .B(n2480), .C(n2501), .D(n2363), .Z(
        n2601) );
  HS65_LS_AOI222X2 U10850 ( .A(n903), .B(n917), .C(n899), .D(n929), .E(n915), 
        .F(n906), .Z(n2598) );
  HS65_LS_NOR4ABX2 U10851 ( .A(n2222), .B(n2223), .C(n2224), .D(n2225), .Z(
        n2148) );
  HS65_LS_NAND4ABX3 U10852 ( .A(n1934), .B(n2057), .C(n2116), .D(n2073), .Z(
        n2224) );
  HS65_LS_NAND4ABX3 U10853 ( .A(n2010), .B(n2104), .C(n2125), .D(n1987), .Z(
        n2225) );
  HS65_LS_AND4X3 U10854 ( .A(n2229), .B(n2004), .C(n2097), .D(n2031), .Z(n2223) );
  HS65_LS_NOR4ABX2 U10855 ( .A(n1470), .B(n1471), .C(n1472), .D(n1473), .Z(
        n1396) );
  HS65_LS_NAND4ABX3 U10856 ( .A(n1258), .B(n1352), .C(n1373), .D(n1235), .Z(
        n1473) );
  HS65_LS_NAND4ABX3 U10857 ( .A(n1182), .B(n1305), .C(n1364), .D(n1321), .Z(
        n1472) );
  HS65_LS_AND4X3 U10858 ( .A(n1477), .B(n1252), .C(n1345), .D(n1279), .Z(n1471) );
  HS65_LS_NOR4ABX2 U10859 ( .A(n4206), .B(n4207), .C(n4208), .D(n4209), .Z(
        n4060) );
  HS65_LS_NAND4ABX3 U10860 ( .A(n3117), .B(n3463), .C(n3533), .D(n3092), .Z(
        n4209) );
  HS65_LS_NAND4ABX3 U10861 ( .A(n2955), .B(n3479), .C(n3458), .D(n3495), .Z(
        n4208) );
  HS65_LS_AOI222X2 U10862 ( .A(n218), .B(n191), .C(n214), .D(n205), .E(n203), 
        .F(n223), .Z(n4206) );
  HS65_LS_NAND2X2 U10863 ( .A(n458), .B(n487), .Z(n5424) );
  HS65_LS_NAND2X2 U10864 ( .A(n239), .B(n268), .Z(n5309) );
  HS65_LS_NAND2X2 U10865 ( .A(n281), .B(n310), .Z(n7016) );
  HS65_LS_NAND2X2 U10866 ( .A(n683), .B(n704), .Z(n5193) );
  HS65_LS_NAND2X2 U10867 ( .A(n60), .B(n89), .Z(n6901) );
  HS65_LS_NAND2X2 U10868 ( .A(n501), .B(n522), .Z(n6785) );
  HS65_LS_NOR3X1 U10869 ( .A(n8269), .B(n8021), .C(n8289), .Z(n8953) );
  HS65_LS_NOR3X1 U10870 ( .A(n8573), .B(n8063), .C(n8593), .Z(n8893) );
  HS65_LS_NAND2X2 U10871 ( .A(n18), .B(n36), .Z(n5045) );
  HS65_LS_NAND2X2 U10872 ( .A(n544), .B(n562), .Z(n6638) );
  HS65_LS_NAND2X2 U10873 ( .A(n55), .B(n85), .Z(n6938) );
  HS65_LS_NAND2X2 U10874 ( .A(n234), .B(n264), .Z(n5346) );
  HS65_LS_NAND2X2 U10875 ( .A(n453), .B(n483), .Z(n5461) );
  HS65_LS_NAND2X2 U10876 ( .A(n276), .B(n306), .Z(n7053) );
  HS65_LS_NAND2X2 U10877 ( .A(n549), .B(n563), .Z(n6717) );
  HS65_LS_NAND2X2 U10878 ( .A(n505), .B(n519), .Z(n6822) );
  HS65_LS_NAND2X2 U10879 ( .A(n23), .B(n37), .Z(n5124) );
  HS65_LS_NAND2X2 U10880 ( .A(n687), .B(n701), .Z(n5230) );
  HS65_LS_NAND2X2 U10881 ( .A(n97), .B(n128), .Z(n7925) );
  HS65_LS_NAND2X2 U10882 ( .A(n584), .B(n615), .Z(n7826) );
  HS65_LS_NAND4ABX3 U10883 ( .A(n4107), .B(n4108), .C(n4109), .D(n4110), .Z(
        n3924) );
  HS65_LS_AOI222X2 U10884 ( .A(n145), .B(n175), .C(n155), .D(n180), .E(n160), 
        .F(n174), .Z(n4109) );
  HS65_LS_NOR4ABX2 U10885 ( .A(n3628), .B(n3656), .C(n3261), .D(n3636), .Z(
        n4110) );
  HS65_LS_NAND4ABX3 U10886 ( .A(n3556), .B(n3246), .C(n4111), .D(n3566), .Z(
        n4108) );
  HS65_LS_NAND4ABX3 U10887 ( .A(n1836), .B(n1837), .C(n1838), .D(n1839), .Z(
        n1764) );
  HS65_LS_NAND4ABX3 U10888 ( .A(n1650), .B(n1603), .C(n1663), .D(n1842), .Z(
        n1837) );
  HS65_LS_AOI222X2 U10889 ( .A(n828), .B(n835), .C(n839), .D(n812), .E(n819), 
        .F(n847), .Z(n1838) );
  HS65_LS_MX41X4 U10890 ( .D0(n848), .S0(n813), .D1(n815), .S1(n843), .D2(n824), .S2(n834), .D3(n845), .S3(n814), .Z(n1836) );
  HS65_LS_NAND4ABX3 U10891 ( .A(n2588), .B(n2589), .C(n2590), .D(n2591), .Z(
        n2516) );
  HS65_LS_NAND4ABX3 U10892 ( .A(n2402), .B(n2355), .C(n2415), .D(n2594), .Z(
        n2589) );
  HS65_LS_AOI222X2 U10893 ( .A(n910), .B(n917), .C(n921), .D(n894), .E(n901), 
        .F(n929), .Z(n2590) );
  HS65_LS_MX41X4 U10894 ( .D0(n930), .S0(n895), .D1(n897), .S1(n925), .D2(n906), .S2(n916), .D3(n927), .S3(n896), .Z(n2588) );
  HS65_LS_NAND4ABX3 U10895 ( .A(n2212), .B(n2213), .C(n2214), .D(n2215), .Z(
        n2140) );
  HS65_LS_NAND4ABX3 U10896 ( .A(n2026), .B(n1979), .C(n2039), .D(n2218), .Z(
        n2213) );
  HS65_LS_AOI222X2 U10897 ( .A(n787), .B(n794), .C(n798), .D(n771), .E(n778), 
        .F(n806), .Z(n2214) );
  HS65_LS_NOR4ABX2 U10898 ( .A(n1997), .B(n2067), .C(n2092), .D(n2085), .Z(
        n2215) );
  HS65_LS_NAND4ABX3 U10899 ( .A(n1460), .B(n1461), .C(n1462), .D(n1463), .Z(
        n1388) );
  HS65_LS_NAND4ABX3 U10900 ( .A(n1274), .B(n1227), .C(n1287), .D(n1466), .Z(
        n1461) );
  HS65_LS_AOI222X2 U10901 ( .A(n869), .B(n876), .C(n880), .D(n853), .E(n860), 
        .F(n888), .Z(n1462) );
  HS65_LS_NOR4ABX2 U10902 ( .A(n1245), .B(n1315), .C(n1340), .D(n1333), .Z(
        n1463) );
  HS65_LS_NAND2X2 U10903 ( .A(n398), .B(n367), .Z(n8116) );
  HS65_LS_NAND2X2 U10904 ( .A(n906), .B(n928), .Z(n2459) );
  HS65_LS_NAND2X2 U10905 ( .A(n824), .B(n846), .Z(n1707) );
  HS65_LS_IVX2 U10906 ( .A(n1128), .Z(n886) );
  HS65_LS_IVX2 U10907 ( .A(n1880), .Z(n804) );
  HS65_LS_IVX2 U10908 ( .A(n2256), .Z(n927) );
  HS65_LS_NAND2X2 U10909 ( .A(n172), .B(n143), .Z(n3595) );
  HS65_LS_IVX2 U10910 ( .A(n1504), .Z(n845) );
  HS65_LS_NAND2X2 U10911 ( .A(n783), .B(n805), .Z(n2083) );
  HS65_LS_NAND2X2 U10912 ( .A(n865), .B(n887), .Z(n1331) );
  HS65_LS_NAND2X2 U10913 ( .A(n91), .B(n63), .Z(n6343) );
  HS65_LS_NAND2X2 U10914 ( .A(n489), .B(n461), .Z(n4789) );
  HS65_LS_NAND2X2 U10915 ( .A(n312), .B(n284), .Z(n6382) );
  HS65_LS_NAND2X2 U10916 ( .A(n270), .B(n242), .Z(n4750) );
  HS65_LS_NAND2X2 U10917 ( .A(n706), .B(n679), .Z(n4643) );
  HS65_LS_NAND2X2 U10918 ( .A(n524), .B(n497), .Z(n6236) );
  HS65_LS_NAND4ABX3 U10919 ( .A(n7261), .B(n7262), .C(n7263), .D(n7264), .Z(
        n7080) );
  HS65_LS_AOI222X2 U10920 ( .A(n536), .B(n555), .C(n550), .D(n564), .E(n548), 
        .F(n557), .Z(n7263) );
  HS65_LS_NAND4ABX3 U10921 ( .A(n6158), .B(n6702), .C(n6625), .D(n6304), .Z(
        n7262) );
  HS65_LS_NAND4ABX3 U10922 ( .A(n6281), .B(n6715), .C(n7265), .D(n6324), .Z(
        n7261) );
  HS65_LS_NAND4ABX3 U10923 ( .A(n5669), .B(n5670), .C(n5671), .D(n5672), .Z(
        n5488) );
  HS65_LS_AOI222X2 U10924 ( .A(n10), .B(n29), .C(n24), .D(n38), .E(n22), .F(
        n31), .Z(n5671) );
  HS65_LS_NAND4ABX3 U10925 ( .A(n4565), .B(n5109), .C(n5032), .D(n4711), .Z(
        n5670) );
  HS65_LS_NAND4ABX3 U10926 ( .A(n4688), .B(n5122), .C(n5673), .D(n4731), .Z(
        n5669) );
  HS65_LS_IVX2 U10927 ( .A(n2765), .Z(n364) );
  HS65_LS_NAND2X2 U10928 ( .A(n160), .B(n180), .Z(n3272) );
  HS65_LS_NAND2X2 U10929 ( .A(n424), .B(n441), .Z(n3818) );
  HS65_LS_NAND2X2 U10930 ( .A(n189), .B(n216), .Z(n3458) );
  HS65_LS_NAND2X2 U10931 ( .A(n458), .B(n481), .Z(n5399) );
  HS65_LS_NAND2X2 U10932 ( .A(n239), .B(n262), .Z(n5284) );
  HS65_LS_NAND2X2 U10933 ( .A(n281), .B(n304), .Z(n6991) );
  HS65_LS_NAND2X2 U10934 ( .A(n683), .B(n700), .Z(n5167) );
  HS65_LS_NAND2X2 U10935 ( .A(n60), .B(n83), .Z(n6876) );
  HS65_LS_NAND2X2 U10936 ( .A(n501), .B(n518), .Z(n6759) );
  HS65_LS_NAND2X2 U10937 ( .A(n920), .B(n903), .Z(n2416) );
  HS65_LS_NAND2X2 U10938 ( .A(n838), .B(n821), .Z(n1664) );
  HS65_LS_NAND2X2 U10939 ( .A(n669), .B(n645), .Z(n3747) );
  HS65_LS_NAND2X2 U10940 ( .A(n879), .B(n862), .Z(n1288) );
  HS65_LS_NAND2X2 U10941 ( .A(n797), .B(n780), .Z(n2040) );
  HS65_LS_IVX2 U10942 ( .A(n2740), .Z(n187) );
  HS65_LS_NAND2X2 U10943 ( .A(n56), .B(n83), .Z(n6937) );
  HS65_LS_NAND2X2 U10944 ( .A(n235), .B(n262), .Z(n5345) );
  HS65_LS_NAND2X2 U10945 ( .A(n454), .B(n481), .Z(n5460) );
  HS65_LS_NAND2X2 U10946 ( .A(n277), .B(n304), .Z(n7052) );
  HS65_LS_NAND2X2 U10947 ( .A(n506), .B(n518), .Z(n6821) );
  HS65_LS_NAND2X2 U10948 ( .A(n688), .B(n700), .Z(n5229) );
  HS65_LS_NAND2X2 U10949 ( .A(n918), .B(n903), .Z(n2458) );
  HS65_LS_NAND2X2 U10950 ( .A(n836), .B(n821), .Z(n1706) );
  HS65_LS_NAND2X2 U10951 ( .A(n68), .B(n85), .Z(n6926) );
  HS65_LS_NAND2X2 U10952 ( .A(n247), .B(n264), .Z(n5334) );
  HS65_LS_NAND2X2 U10953 ( .A(n466), .B(n483), .Z(n5449) );
  HS65_LS_NAND2X2 U10954 ( .A(n289), .B(n306), .Z(n7041) );
  HS65_LS_NAND2X2 U10955 ( .A(n536), .B(n563), .Z(n6689) );
  HS65_LS_NAND2X2 U10956 ( .A(n493), .B(n519), .Z(n6810) );
  HS65_LS_NAND2X2 U10957 ( .A(n10), .B(n37), .Z(n5096) );
  HS65_LS_NAND2X2 U10958 ( .A(n675), .B(n701), .Z(n5218) );
  HS65_LS_NAND2X2 U10959 ( .A(n154), .B(n167), .Z(n3048) );
  HS65_LS_NAND2X2 U10960 ( .A(n877), .B(n862), .Z(n1330) );
  HS65_LS_NAND2X2 U10961 ( .A(n795), .B(n780), .Z(n2082) );
  HS65_LS_NAND2X2 U10962 ( .A(n833), .B(n821), .Z(n1637) );
  HS65_LS_NAND2X2 U10963 ( .A(n915), .B(n903), .Z(n2389) );
  HS65_LS_NAND4ABX3 U10964 ( .A(n4253), .B(n4254), .C(n4255), .D(n4256), .Z(
        n2890) );
  HS65_LS_NAND4ABX3 U10965 ( .A(n3336), .B(n3159), .C(n3722), .D(n3701), .Z(
        n4254) );
  HS65_LS_NOR4ABX2 U10966 ( .A(n3764), .B(n3708), .C(n3327), .D(n3745), .Z(
        n4256) );
  HS65_LS_AOI222X2 U10967 ( .A(n649), .B(n656), .C(n671), .D(n641), .E(n650), 
        .F(n655), .Z(n4255) );
  HS65_LS_NAND2X2 U10968 ( .A(n329), .B(n344), .Z(n8616) );
  HS65_LS_NAND2X2 U10969 ( .A(n550), .B(n562), .Z(n6716) );
  HS65_LS_NAND2X2 U10970 ( .A(n24), .B(n36), .Z(n5123) );
  HS65_LS_NAND2X2 U10971 ( .A(n874), .B(n862), .Z(n1261) );
  HS65_LS_NAND2X2 U10972 ( .A(n792), .B(n780), .Z(n2013) );
  HS65_LS_NAND2X2 U10973 ( .A(n568), .B(n540), .Z(n6159) );
  HS65_LS_NAND2X2 U10974 ( .A(n42), .B(n14), .Z(n4566) );
  HS65_LS_NAND2X2 U10975 ( .A(n910), .B(n924), .Z(n2483) );
  HS65_LS_NAND2X2 U10976 ( .A(n828), .B(n842), .Z(n1731) );
  HS65_LS_NAND4ABX3 U10977 ( .A(n2426), .B(n2427), .C(n2428), .D(n2429), .Z(
        n2316) );
  HS65_LS_NOR3AX2 U10978 ( .A(n2434), .B(n2435), .C(n2436), .Z(n2428) );
  HS65_LS_NAND4ABX3 U10979 ( .A(n2441), .B(n2442), .C(n2443), .D(n2444), .Z(
        n2426) );
  HS65_LS_NOR4ABX2 U10980 ( .A(n2430), .B(n2431), .C(n2432), .D(n2433), .Z(
        n2429) );
  HS65_LS_NAND4ABX3 U10981 ( .A(n1674), .B(n1675), .C(n1676), .D(n1677), .Z(
        n1564) );
  HS65_LS_NOR3AX2 U10982 ( .A(n1682), .B(n1683), .C(n1684), .Z(n1676) );
  HS65_LS_NAND4ABX3 U10983 ( .A(n1689), .B(n1690), .C(n1691), .D(n1692), .Z(
        n1674) );
  HS65_LS_NOR4ABX2 U10984 ( .A(n1678), .B(n1679), .C(n1680), .D(n1681), .Z(
        n1677) );
  HS65_LS_NAND4ABX3 U10985 ( .A(n1298), .B(n1299), .C(n1300), .D(n1301), .Z(
        n1188) );
  HS65_LS_NOR3AX2 U10986 ( .A(n1306), .B(n1307), .C(n1308), .Z(n1300) );
  HS65_LS_NOR4ABX2 U10987 ( .A(n1302), .B(n1303), .C(n1304), .D(n1305), .Z(
        n1301) );
  HS65_LS_NAND4ABX3 U10988 ( .A(n1313), .B(n1314), .C(n1315), .D(n1316), .Z(
        n1298) );
  HS65_LS_NAND4ABX3 U10989 ( .A(n2050), .B(n2051), .C(n2052), .D(n2053), .Z(
        n1940) );
  HS65_LS_NOR3AX2 U10990 ( .A(n2058), .B(n2059), .C(n2060), .Z(n2052) );
  HS65_LS_NOR4ABX2 U10991 ( .A(n2054), .B(n2055), .C(n2056), .D(n2057), .Z(
        n2053) );
  HS65_LS_NAND4ABX3 U10992 ( .A(n2065), .B(n2066), .C(n2067), .D(n2068), .Z(
        n2050) );
  HS65_LS_NAND2X2 U10993 ( .A(n869), .B(n883), .Z(n1355) );
  HS65_LS_NAND2X2 U10994 ( .A(n787), .B(n801), .Z(n2107) );
  HS65_LS_NAND2X2 U10995 ( .A(n440), .B(n419), .Z(n3399) );
  HS65_LS_NAND2X2 U10996 ( .A(n923), .B(n900), .Z(n2492) );
  HS65_LS_NAND2X2 U10997 ( .A(n841), .B(n818), .Z(n1740) );
  HS65_LS_NAND2X2 U10998 ( .A(n882), .B(n859), .Z(n1364) );
  HS65_LS_NAND2X2 U10999 ( .A(n107), .B(n128), .Z(n7918) );
  HS65_LS_NAND2X2 U11000 ( .A(n594), .B(n615), .Z(n7819) );
  HS65_LS_NAND4ABX3 U11001 ( .A(n7449), .B(n7450), .C(n7451), .D(n7452), .Z(
        n7139) );
  HS65_LS_AOI222X2 U11002 ( .A(n68), .B(n81), .C(n56), .D(n84), .E(n62), .F(
        n82), .Z(n7451) );
  HS65_LS_NAND4ABX3 U11003 ( .A(n6342), .B(n6952), .C(n6862), .D(n6520), .Z(
        n7450) );
  HS65_LS_NAND4ABX3 U11004 ( .A(n6499), .B(n6936), .C(n7455), .D(n6538), .Z(
        n7449) );
  HS65_LS_NAND4ABX3 U11005 ( .A(n5916), .B(n5917), .C(n5918), .D(n5919), .Z(
        n5568) );
  HS65_LS_AOI222X2 U11006 ( .A(n466), .B(n479), .C(n454), .D(n482), .E(n460), 
        .F(n480), .Z(n5918) );
  HS65_LS_NAND4ABX3 U11007 ( .A(n4788), .B(n5475), .C(n5385), .D(n4981), .Z(
        n5917) );
  HS65_LS_NAND4ABX3 U11008 ( .A(n4960), .B(n5459), .C(n5922), .D(n4999), .Z(
        n5916) );
  HS65_LS_NAND4ABX3 U11009 ( .A(n7508), .B(n7509), .C(n7510), .D(n7511), .Z(
        n7160) );
  HS65_LS_AOI222X2 U11010 ( .A(n289), .B(n302), .C(n277), .D(n305), .E(n283), 
        .F(n303), .Z(n7510) );
  HS65_LS_NAND4ABX3 U11011 ( .A(n6381), .B(n7067), .C(n6977), .D(n6574), .Z(
        n7509) );
  HS65_LS_NAND4ABX3 U11012 ( .A(n6553), .B(n7051), .C(n7514), .D(n6592), .Z(
        n7508) );
  HS65_LS_NAND4ABX3 U11013 ( .A(n5857), .B(n5858), .C(n5859), .D(n5860), .Z(
        n5547) );
  HS65_LS_AOI222X2 U11014 ( .A(n247), .B(n260), .C(n235), .D(n263), .E(n241), 
        .F(n261), .Z(n5859) );
  HS65_LS_NAND4ABX3 U11015 ( .A(n4749), .B(n5360), .C(n5270), .D(n4927), .Z(
        n5858) );
  HS65_LS_NAND4ABX3 U11016 ( .A(n4906), .B(n5344), .C(n5863), .D(n4945), .Z(
        n5857) );
  HS65_LS_NAND4ABX3 U11017 ( .A(n5699), .B(n5700), .C(n5701), .D(n5702), .Z(
        n5504) );
  HS65_LS_AOI222X2 U11018 ( .A(n675), .B(n693), .C(n688), .D(n702), .E(n686), 
        .F(n695), .Z(n5701) );
  HS65_LS_NAND4ABX3 U11019 ( .A(n4642), .B(n5245), .C(n5153), .D(n4851), .Z(
        n5700) );
  HS65_LS_NAND4ABX3 U11020 ( .A(n4829), .B(n5228), .C(n5703), .D(n4871), .Z(
        n5699) );
  HS65_LS_NAND4ABX3 U11021 ( .A(n7291), .B(n7292), .C(n7293), .D(n7294), .Z(
        n7096) );
  HS65_LS_AOI222X2 U11022 ( .A(n493), .B(n511), .C(n506), .D(n520), .E(n504), 
        .F(n513), .Z(n7293) );
  HS65_LS_NAND4ABX3 U11023 ( .A(n6235), .B(n6837), .C(n6745), .D(n6444), .Z(
        n7292) );
  HS65_LS_NAND4ABX3 U11024 ( .A(n6422), .B(n6820), .C(n7295), .D(n6464), .Z(
        n7291) );
  HS65_LS_NAND2X2 U11025 ( .A(n800), .B(n777), .Z(n2116) );
  HS65_LS_NAND2X2 U11026 ( .A(n543), .B(n558), .Z(n6712) );
  HS65_LS_NAND2X2 U11027 ( .A(n17), .B(n32), .Z(n5119) );
  HS65_LS_NOR4ABX2 U11028 ( .A(n2275), .B(n2276), .C(n2277), .D(n2278), .Z(
        n2274) );
  HS65_LS_AOI212X2 U11029 ( .A(n918), .B(n899), .C(n930), .D(n908), .E(n2279), 
        .Z(n2276) );
  HS65_LS_NOR4ABX2 U11030 ( .A(n1523), .B(n1524), .C(n1525), .D(n1526), .Z(
        n1522) );
  HS65_LS_AOI212X2 U11031 ( .A(n836), .B(n817), .C(n848), .D(n826), .E(n1527), 
        .Z(n1524) );
  HS65_LS_NOR4ABX2 U11032 ( .A(n1147), .B(n1148), .C(n1149), .D(n1150), .Z(
        n1146) );
  HS65_LS_AOI212X2 U11033 ( .A(n877), .B(n858), .C(n889), .D(n867), .E(n1151), 
        .Z(n1148) );
  HS65_LS_NOR4ABX2 U11034 ( .A(n1899), .B(n1900), .C(n1901), .D(n1902), .Z(
        n1898) );
  HS65_LS_AOI212X2 U11035 ( .A(n795), .B(n776), .C(n807), .D(n785), .E(n1903), 
        .Z(n1900) );
  HS65_LS_NAND2X2 U11036 ( .A(n193), .B(n218), .Z(n3444) );
  HS65_LS_NAND4ABX3 U11037 ( .A(n4312), .B(n4313), .C(n4314), .D(n4315), .Z(
        n2845) );
  HS65_LS_AOI222X2 U11038 ( .A(n425), .B(n432), .C(n447), .D(n417), .E(n426), 
        .F(n431), .Z(n4314) );
  HS65_LS_NOR4ABX2 U11039 ( .A(n3881), .B(n3388), .C(n3824), .D(n3862), .Z(
        n4315) );
  HS65_LS_NAND4ABX3 U11040 ( .A(n3839), .B(n3200), .C(n3399), .D(n3817), .Z(
        n4313) );
  HS65_LS_NAND2X2 U11041 ( .A(n194), .B(n218), .Z(n3505) );
  HS65_LS_NAND2X2 U11042 ( .A(n65), .B(n79), .Z(n6933) );
  HS65_LS_NAND2X2 U11043 ( .A(n244), .B(n258), .Z(n5341) );
  HS65_LS_NAND2X2 U11044 ( .A(n463), .B(n477), .Z(n5456) );
  HS65_LS_NAND2X2 U11045 ( .A(n286), .B(n300), .Z(n7048) );
  HS65_LS_NAND2X2 U11046 ( .A(n500), .B(n514), .Z(n6817) );
  HS65_LS_NAND2X2 U11047 ( .A(n682), .B(n696), .Z(n5225) );
  HS65_LS_NAND4ABX3 U11048 ( .A(n1825), .B(n1826), .C(n1827), .D(n1828), .Z(
        n1501) );
  HS65_LS_AOI222X2 U11049 ( .A(n835), .B(n812), .C(n815), .D(n839), .E(n848), 
        .F(n826), .Z(n1827) );
  HS65_LS_NAND4ABX3 U11050 ( .A(n1626), .B(n1560), .C(n1682), .D(n1739), .Z(
        n1826) );
  HS65_LS_NOR4ABX2 U11051 ( .A(n1724), .B(n1616), .C(n1729), .D(n1705), .Z(
        n1828) );
  HS65_LS_NAND4ABX3 U11052 ( .A(n2577), .B(n2578), .C(n2579), .D(n2580), .Z(
        n2253) );
  HS65_LS_AOI222X2 U11053 ( .A(n917), .B(n894), .C(n897), .D(n921), .E(n930), 
        .F(n908), .Z(n2579) );
  HS65_LS_NAND4ABX3 U11054 ( .A(n2378), .B(n2312), .C(n2434), .D(n2491), .Z(
        n2578) );
  HS65_LS_NOR4ABX2 U11055 ( .A(n2476), .B(n2368), .C(n2481), .D(n2457), .Z(
        n2580) );
  HS65_LS_NAND4ABX3 U11056 ( .A(n1449), .B(n1450), .C(n1451), .D(n1452), .Z(
        n1125) );
  HS65_LS_AOI222X2 U11057 ( .A(n876), .B(n853), .C(n856), .D(n880), .E(n889), 
        .F(n867), .Z(n1451) );
  HS65_LS_NAND4ABX3 U11058 ( .A(n1250), .B(n1184), .C(n1306), .D(n1363), .Z(
        n1450) );
  HS65_LS_NOR4ABX2 U11059 ( .A(n1348), .B(n1240), .C(n1353), .D(n1329), .Z(
        n1452) );
  HS65_LS_NAND4ABX3 U11060 ( .A(n2201), .B(n2202), .C(n2203), .D(n2204), .Z(
        n1877) );
  HS65_LS_AOI222X2 U11061 ( .A(n794), .B(n771), .C(n774), .D(n798), .E(n807), 
        .F(n785), .Z(n2203) );
  HS65_LS_NAND4ABX3 U11062 ( .A(n2002), .B(n1936), .C(n2058), .D(n2115), .Z(
        n2202) );
  HS65_LS_NOR4ABX2 U11063 ( .A(n2100), .B(n1992), .C(n2105), .D(n2081), .Z(
        n2204) );
  HS65_LS_NAND2X2 U11064 ( .A(n203), .B(n218), .Z(n3120) );
  HS65_LS_IVX2 U11065 ( .A(n2763), .Z(n362) );
  HS65_LS_NAND4ABX3 U11066 ( .A(n4129), .B(n4130), .C(n4131), .D(n4132), .Z(
        n4098) );
  HS65_LS_NAND4ABX3 U11067 ( .A(n3572), .B(n3579), .C(n3594), .D(n4133), .Z(
        n4129) );
  HS65_LS_NAND4ABX3 U11068 ( .A(n3271), .B(n3284), .C(n3258), .D(n3035), .Z(
        n4130) );
  HS65_LS_AOI222X2 U11069 ( .A(n145), .B(n180), .C(n177), .D(n155), .E(n182), 
        .F(n144), .Z(n4131) );
  HS65_LS_IVX2 U11070 ( .A(n2832), .Z(n452) );
  HS65_LS_IVX2 U11071 ( .A(n2824), .Z(n275) );
  HS65_LS_NAND2X2 U11072 ( .A(n330), .B(n350), .Z(n8375) );
  HS65_LS_IVX2 U11073 ( .A(n2652), .Z(n186) );
  HS65_LS_NOR4ABX2 U11074 ( .A(n1765), .B(n1787), .C(n1502), .D(n1788), .Z(
        n1786) );
  HS65_LS_AOI212X2 U11075 ( .A(n848), .B(n821), .C(n815), .D(n841), .E(n1773), 
        .Z(n1787) );
  HS65_LS_NOR4ABX2 U11076 ( .A(n2517), .B(n2539), .C(n2254), .D(n2540), .Z(
        n2538) );
  HS65_LS_AOI212X2 U11077 ( .A(n930), .B(n903), .C(n897), .D(n923), .E(n2525), 
        .Z(n2539) );
  HS65_LS_NOR4ABX2 U11078 ( .A(n1389), .B(n1411), .C(n1126), .D(n1412), .Z(
        n1410) );
  HS65_LS_AOI212X2 U11079 ( .A(n889), .B(n862), .C(n856), .D(n882), .E(n1397), 
        .Z(n1411) );
  HS65_LS_NOR4ABX2 U11080 ( .A(n2141), .B(n2163), .C(n1878), .D(n2164), .Z(
        n2162) );
  HS65_LS_AOI212X2 U11081 ( .A(n807), .B(n780), .C(n774), .D(n800), .E(n2149), 
        .Z(n2163) );
  HS65_LS_NOR4ABX2 U11082 ( .A(n3925), .B(n3994), .C(n3995), .D(n3996), .Z(
        n3993) );
  HS65_LS_AOI212X2 U11083 ( .A(n171), .B(n144), .C(n143), .D(n177), .E(n3997), 
        .Z(n3994) );
  HS65_LS_NOR4ABX2 U11084 ( .A(n3907), .B(n3932), .C(n3933), .D(n3934), .Z(
        n3931) );
  HS65_LS_AOI212X2 U11085 ( .A(n190), .B(n218), .C(n222), .D(n189), .E(n3935), 
        .Z(n3932) );
  HS65_LS_NAND2X2 U11086 ( .A(n160), .B(n176), .Z(n3643) );
  HS65_LS_NAND2X2 U11087 ( .A(n21), .B(n32), .Z(n4691) );
  HS65_LS_NAND2X2 U11088 ( .A(n547), .B(n558), .Z(n6284) );
  HS65_LS_NAND2X2 U11089 ( .A(n645), .B(n659), .Z(n3773) );
  HS65_LS_NAND2X2 U11090 ( .A(n156), .B(n172), .Z(n3570) );
  HS65_LS_NAND2X2 U11091 ( .A(n147), .B(n177), .Z(n3594) );
  HS65_LS_NAND2X2 U11092 ( .A(n671), .B(n647), .Z(n3701) );
  HS65_LS_NAND2X2 U11093 ( .A(n61), .B(n79), .Z(n6501) );
  HS65_LS_NAND2X2 U11094 ( .A(n282), .B(n300), .Z(n6555) );
  HS65_LS_NAND2X2 U11095 ( .A(n240), .B(n258), .Z(n4908) );
  HS65_LS_NAND2X2 U11096 ( .A(n459), .B(n477), .Z(n4962) );
  HS65_LS_NAND2X2 U11097 ( .A(n685), .B(n696), .Z(n4831) );
  HS65_LS_NAND2X2 U11098 ( .A(n503), .B(n514), .Z(n6424) );
  HS65_LS_NOR2X2 U11099 ( .A(n900), .B(n895), .Z(n2287) );
  HS65_LS_NOR2X2 U11100 ( .A(n818), .B(n813), .Z(n1535) );
  HS65_LS_NOR2X2 U11101 ( .A(n859), .B(n854), .Z(n1159) );
  HS65_LS_NOR2X2 U11102 ( .A(n777), .B(n772), .Z(n1911) );
  HS65_LS_NAND2X2 U11103 ( .A(n195), .B(n213), .Z(n3533) );
  HS65_LS_NAND2X2 U11104 ( .A(n419), .B(n439), .Z(n3805) );
  HS65_LS_NAND2X2 U11105 ( .A(n846), .B(n822), .Z(n1749) );
  HS65_LS_NAND2X2 U11106 ( .A(n928), .B(n904), .Z(n2501) );
  HS65_LS_NAND2X2 U11107 ( .A(n887), .B(n863), .Z(n1373) );
  HS65_LS_NAND2X2 U11108 ( .A(n805), .B(n781), .Z(n2125) );
  HS65_LS_NAND2X2 U11109 ( .A(n422), .B(n439), .Z(n3863) );
  HS65_LS_NAND2X2 U11110 ( .A(n410), .B(n439), .Z(n3409) );
  HS65_LS_NAND2X2 U11111 ( .A(n421), .B(n435), .Z(n3890) );
  HS65_LS_NAND2X2 U11112 ( .A(n159), .B(n175), .Z(n3266) );
  HS65_LS_NOR4ABX2 U11113 ( .A(n7688), .B(n7689), .C(n7690), .D(n7631), .Z(
        n7678) );
  HS65_LS_NOR4ABX2 U11114 ( .A(n7726), .B(n7727), .C(n7728), .D(n7659), .Z(
        n7716) );
  HS65_LS_IVX2 U11115 ( .A(n2757), .Z(n629) );
  HS65_LS_NAND2X2 U11116 ( .A(n40), .B(n18), .Z(n5071) );
  HS65_LS_NAND2X2 U11117 ( .A(n566), .B(n544), .Z(n6664) );
  HS65_LS_NAND2X2 U11118 ( .A(n343), .B(n336), .Z(n8539) );
  HS65_LS_NAND2X2 U11119 ( .A(n376), .B(n399), .Z(n8091) );
  HS65_LS_NAND2X2 U11120 ( .A(n370), .B(n399), .Z(n8239) );
  HS65_LS_IVX2 U11121 ( .A(n2645), .Z(n188) );
  HS65_LS_NOR4ABX2 U11122 ( .A(n5627), .B(n5561), .C(n4507), .D(n5556), .Z(
        n5890) );
  HS65_LS_NOR4ABX2 U11123 ( .A(n5600), .B(n5540), .C(n4461), .D(n5535), .Z(
        n5831) );
  HS65_LS_NOR4ABX2 U11124 ( .A(n5583), .B(n5684), .C(n5685), .D(n5502), .Z(
        n5680) );
  HS65_LS_NOR4ABX2 U11125 ( .A(n7219), .B(n7153), .C(n6100), .D(n7148), .Z(
        n7482) );
  HS65_LS_NOR4ABX2 U11126 ( .A(n7192), .B(n7132), .C(n6054), .D(n7127), .Z(
        n7423) );
  HS65_LS_NOR4ABX2 U11127 ( .A(n7175), .B(n7276), .C(n7277), .D(n7094), .Z(
        n7272) );
  HS65_LS_NOR4ABX2 U11128 ( .A(n7780), .B(n7781), .C(n7782), .D(n7783), .Z(
        n7769) );
  HS65_LS_NAND2X2 U11129 ( .A(n402), .B(n373), .Z(n8312) );
  HS65_LS_IVX2 U11130 ( .A(n2790), .Z(n579) );
  HS65_LS_NOR4ABX2 U11131 ( .A(n2978), .B(n2979), .C(n2980), .D(n2981), .Z(
        n2977) );
  HS65_LS_AO212X4 U11132 ( .A(n646), .B(n660), .C(n650), .D(n655), .E(n2982), 
        .Z(n2980) );
  HS65_LS_NOR4ABX2 U11133 ( .A(n2866), .B(n2867), .C(n2868), .D(n2869), .Z(
        n2865) );
  HS65_LS_AO212X4 U11134 ( .A(n194), .B(n214), .C(n190), .D(n228), .E(n2870), 
        .Z(n2868) );
  HS65_LS_NOR4ABX2 U11135 ( .A(n2996), .B(n2997), .C(n2998), .D(n2999), .Z(
        n2995) );
  HS65_LS_AO212X4 U11136 ( .A(n422), .B(n436), .C(n426), .D(n431), .E(n3000), 
        .Z(n2998) );
  HS65_LS_NAND4ABX3 U11137 ( .A(n6639), .B(n6640), .C(n6641), .D(n6642), .Z(
        n6299) );
  HS65_LS_OR4X4 U11138 ( .A(n6655), .B(n6656), .C(n6657), .D(n6658), .Z(n6639)
         );
  HS65_LS_NAND3X2 U11139 ( .A(n6651), .B(n6652), .C(n6653), .Z(n6640) );
  HS65_LS_NOR4ABX2 U11140 ( .A(n6643), .B(n6644), .C(n545), .D(n6645), .Z(
        n6642) );
  HS65_LS_NAND4ABX3 U11141 ( .A(n5046), .B(n5047), .C(n5048), .D(n5049), .Z(
        n4706) );
  HS65_LS_OR4X4 U11142 ( .A(n5062), .B(n5063), .C(n5064), .D(n5065), .Z(n5046)
         );
  HS65_LS_NAND3X2 U11143 ( .A(n5058), .B(n5059), .C(n5060), .Z(n5047) );
  HS65_LS_NOR4ABX2 U11144 ( .A(n5050), .B(n5051), .C(n19), .D(n5052), .Z(n5049) );
  HS65_LS_NAND4ABX3 U11145 ( .A(n3368), .B(n3369), .C(n3370), .D(n3371), .Z(
        n3182) );
  HS65_LS_NAND4ABX3 U11146 ( .A(n3397), .B(n3398), .C(n3399), .D(n3400), .Z(
        n3369) );
  HS65_LS_NOR4ABX2 U11147 ( .A(n3372), .B(n3373), .C(n3374), .D(n3375), .Z(
        n3371) );
  HS65_LS_MX41X4 U11148 ( .D0(n423), .S0(n441), .D1(n426), .S1(n447), .D2(n410), .S2(n434), .D3(n415), .S3(n443), .Z(n3368) );
  HS65_LS_NAND4ABX3 U11149 ( .A(n6877), .B(n6878), .C(n6879), .D(n6880), .Z(
        n6515) );
  HS65_LS_OR4X4 U11150 ( .A(n6892), .B(n6893), .C(n6894), .D(n6895), .Z(n6877)
         );
  HS65_LS_NOR4ABX2 U11151 ( .A(n6881), .B(n6882), .C(n6883), .D(n6884), .Z(
        n6880) );
  HS65_LS_NAND3X2 U11152 ( .A(n6889), .B(n6890), .C(n6891), .Z(n6878) );
  HS65_LS_NAND4ABX3 U11153 ( .A(n5285), .B(n5286), .C(n5287), .D(n5288), .Z(
        n4922) );
  HS65_LS_OR4X4 U11154 ( .A(n5300), .B(n5301), .C(n5302), .D(n5303), .Z(n5285)
         );
  HS65_LS_NOR4ABX2 U11155 ( .A(n5289), .B(n5290), .C(n5291), .D(n5292), .Z(
        n5288) );
  HS65_LS_NAND3X2 U11156 ( .A(n5297), .B(n5298), .C(n5299), .Z(n5286) );
  HS65_LS_NAND4ABX3 U11157 ( .A(n5400), .B(n5401), .C(n5402), .D(n5403), .Z(
        n4976) );
  HS65_LS_OR4X4 U11158 ( .A(n5415), .B(n5416), .C(n5417), .D(n5418), .Z(n5400)
         );
  HS65_LS_NOR4ABX2 U11159 ( .A(n5404), .B(n5405), .C(n5406), .D(n5407), .Z(
        n5403) );
  HS65_LS_NAND3X2 U11160 ( .A(n5412), .B(n5413), .C(n5414), .Z(n5401) );
  HS65_LS_NAND4ABX3 U11161 ( .A(n6992), .B(n6993), .C(n6994), .D(n6995), .Z(
        n6569) );
  HS65_LS_OR4X4 U11162 ( .A(n7007), .B(n7008), .C(n7009), .D(n7010), .Z(n6992)
         );
  HS65_LS_NOR4ABX2 U11163 ( .A(n6996), .B(n6997), .C(n6998), .D(n6999), .Z(
        n6995) );
  HS65_LS_NAND3X2 U11164 ( .A(n7004), .B(n7005), .C(n7006), .Z(n6993) );
  HS65_LS_NAND4ABX3 U11165 ( .A(n5168), .B(n5169), .C(n5170), .D(n5171), .Z(
        n4846) );
  HS65_LS_OR4X4 U11166 ( .A(n5184), .B(n5185), .C(n5186), .D(n5187), .Z(n5168)
         );
  HS65_LS_NOR4ABX2 U11167 ( .A(n5172), .B(n5173), .C(n5174), .D(n5175), .Z(
        n5171) );
  HS65_LS_NAND3X2 U11168 ( .A(n5180), .B(n5181), .C(n5182), .Z(n5169) );
  HS65_LS_NAND4ABX3 U11169 ( .A(n6760), .B(n6761), .C(n6762), .D(n6763), .Z(
        n6439) );
  HS65_LS_OR4X4 U11170 ( .A(n6776), .B(n6777), .C(n6778), .D(n6779), .Z(n6760)
         );
  HS65_LS_NOR4ABX2 U11171 ( .A(n6764), .B(n6765), .C(n6766), .D(n6767), .Z(
        n6763) );
  HS65_LS_NAND3X2 U11172 ( .A(n6772), .B(n6773), .C(n6774), .Z(n6761) );
  HS65_LS_NAND2X2 U11173 ( .A(n647), .B(n658), .Z(n3750) );
  HS65_LS_IVX2 U11174 ( .A(n2736), .Z(n631) );
  HS65_LS_NAND4ABX3 U11175 ( .A(n3306), .B(n3307), .C(n3308), .D(n3309), .Z(
        n3141) );
  HS65_LS_NAND4ABX3 U11176 ( .A(n3335), .B(n3336), .C(n3337), .D(n3338), .Z(
        n3307) );
  HS65_LS_MX41X4 U11177 ( .D0(n647), .S0(n665), .D1(n650), .S1(n671), .D2(n633), .S2(n658), .D3(n639), .S3(n667), .Z(n3306) );
  HS65_LS_NOR4ABX2 U11178 ( .A(n3310), .B(n3311), .C(n3312), .D(n3313), .Z(
        n3309) );
  HS65_LS_NAND2X2 U11179 ( .A(n837), .B(n823), .Z(n1710) );
  HS65_LS_NAND2X2 U11180 ( .A(n919), .B(n905), .Z(n2462) );
  HS65_LS_IVX2 U11181 ( .A(n2803), .Z(n233) );
  HS65_LS_IVX2 U11182 ( .A(n2795), .Z(n53) );
  HS65_LS_IVX2 U11183 ( .A(n2787), .Z(n577) );
  HS65_LS_NAND2X2 U11184 ( .A(n796), .B(n782), .Z(n2086) );
  HS65_LS_NAND2X2 U11185 ( .A(n878), .B(n864), .Z(n1334) );
  HS65_LS_NAND4ABX3 U11186 ( .A(n3077), .B(n3078), .C(n3079), .D(n3080), .Z(
        n2938) );
  HS65_LS_NAND4ABX3 U11187 ( .A(n3108), .B(n3109), .C(n3110), .D(n3111), .Z(
        n3078) );
  HS65_LS_MX41X4 U11188 ( .D0(n192), .S0(n216), .D1(n190), .S1(n222), .D2(n203), .S2(n225), .D3(n199), .S3(n219), .Z(n3077) );
  HS65_LS_NOR4ABX2 U11189 ( .A(n3081), .B(n3082), .C(n3083), .D(n3084), .Z(
        n3080) );
  HS65_LS_NAND2X2 U11190 ( .A(n897), .B(n919), .Z(n2491) );
  HS65_LS_NAND2X2 U11191 ( .A(n815), .B(n837), .Z(n1739) );
  HS65_LS_NAND2X2 U11192 ( .A(n423), .B(n434), .Z(n3867) );
  HS65_LS_NOR4ABX2 U11193 ( .A(n8082), .B(n7873), .C(n8106), .D(n8012), .Z(
        n8206) );
  HS65_LS_NAND4ABX3 U11194 ( .A(n8575), .B(n8576), .C(n8577), .D(n8578), .Z(
        n8348) );
  HS65_LS_NOR4ABX2 U11195 ( .A(n8583), .B(n8584), .C(n8585), .D(n8586), .Z(
        n8577) );
  HS65_LS_OR4X4 U11196 ( .A(n8590), .B(n8591), .C(n8592), .D(n8593), .Z(n8575)
         );
  HS65_LS_NAND3AX3 U11197 ( .A(n7773), .B(n8587), .C(n8588), .Z(n8576) );
  HS65_LS_NAND2X2 U11198 ( .A(n856), .B(n878), .Z(n1363) );
  HS65_LS_NAND2X2 U11199 ( .A(n774), .B(n796), .Z(n2115) );
  HS65_LS_NAND4ABX3 U11200 ( .A(n8097), .B(n8098), .C(n8099), .D(n8100), .Z(
        n8013) );
  HS65_LS_NAND4ABX3 U11201 ( .A(n8125), .B(n8126), .C(n8127), .D(n8128), .Z(
        n8098) );
  HS65_LS_NOR4ABX2 U11202 ( .A(n8101), .B(n8102), .C(n8103), .D(n8104), .Z(
        n8100) );
  HS65_LS_MX41X4 U11203 ( .D0(n365), .S0(n396), .D1(n395), .S1(n366), .D2(n376), .S2(n388), .D3(n393), .S3(n378), .Z(n8097) );
  HS65_LS_NAND2X2 U11204 ( .A(n222), .B(n192), .Z(n3457) );
  HS65_LS_NOR4ABX2 U11205 ( .A(n2916), .B(n2917), .C(n2918), .D(n2919), .Z(
        n2915) );
  HS65_LS_AO212X4 U11206 ( .A(n149), .B(n168), .C(n182), .D(n144), .E(n2920), 
        .Z(n2918) );
  HS65_LS_NAND4ABX3 U11207 ( .A(n3239), .B(n3240), .C(n3241), .D(n3242), .Z(
        n3030) );
  HS65_LS_NAND4ABX3 U11208 ( .A(n3270), .B(n3271), .C(n3272), .D(n3273), .Z(
        n3240) );
  HS65_LS_NOR4ABX2 U11209 ( .A(n3243), .B(n3244), .C(n3245), .D(n3246), .Z(
        n3242) );
  HS65_LS_MX41X4 U11210 ( .D0(n170), .S0(n147), .D1(n177), .S1(n144), .D2(n158), .S2(n179), .D3(n154), .S3(n174), .Z(n3239) );
  HS65_LS_NOR4ABX2 U11211 ( .A(n7688), .B(n7628), .C(n9009), .D(n7810), .Z(
        n9008) );
  HS65_LS_AO212X4 U11212 ( .A(n608), .B(n585), .C(n592), .D(n611), .E(n7701), 
        .Z(n9009) );
  HS65_LS_NOR4ABX2 U11213 ( .A(n7726), .B(n7656), .C(n9067), .D(n7910), .Z(
        n9066) );
  HS65_LS_AO212X4 U11214 ( .A(n121), .B(n98), .C(n105), .D(n124), .E(n7739), 
        .Z(n9067) );
  HS65_LS_NOR4ABX2 U11215 ( .A(n5554), .B(n5555), .C(n5556), .D(n4506), .Z(
        n5553) );
  HS65_LS_AOI212X2 U11216 ( .A(n474), .B(n461), .C(n468), .D(n471), .E(n5568), 
        .Z(n5555) );
  HS65_LS_NOR4ABX2 U11217 ( .A(n7146), .B(n7147), .C(n7148), .D(n6099), .Z(
        n7145) );
  HS65_LS_AOI212X2 U11218 ( .A(n297), .B(n284), .C(n291), .D(n294), .E(n7160), 
        .Z(n7147) );
  HS65_LS_NOR4ABX2 U11219 ( .A(n7125), .B(n7126), .C(n7127), .D(n6053), .Z(
        n7124) );
  HS65_LS_AOI212X2 U11220 ( .A(n76), .B(n63), .C(n70), .D(n73), .E(n7139), .Z(
        n7126) );
  HS65_LS_NOR4ABX2 U11221 ( .A(n5533), .B(n5534), .C(n5535), .D(n4460), .Z(
        n5532) );
  HS65_LS_AOI212X2 U11222 ( .A(n255), .B(n242), .C(n249), .D(n252), .E(n5547), 
        .Z(n5534) );
  HS65_LS_NOR4ABX2 U11223 ( .A(n7092), .B(n7093), .C(n7094), .D(n7095), .Z(
        n7091) );
  HS65_LS_AOI212X2 U11224 ( .A(n528), .B(n497), .C(n494), .D(n529), .E(n7096), 
        .Z(n7093) );
  HS65_LS_NOR4ABX2 U11225 ( .A(n5484), .B(n5485), .C(n5486), .D(n5487), .Z(
        n5483) );
  HS65_LS_AOI212X2 U11226 ( .A(n46), .B(n14), .C(n11), .D(n47), .E(n5488), .Z(
        n5485) );
  HS65_LS_NOR4ABX2 U11227 ( .A(n7076), .B(n7077), .C(n7078), .D(n7079), .Z(
        n7075) );
  HS65_LS_AOI212X2 U11228 ( .A(n572), .B(n540), .C(n537), .D(n573), .E(n7080), 
        .Z(n7077) );
  HS65_LS_NOR4ABX2 U11229 ( .A(n5500), .B(n5501), .C(n5502), .D(n5503), .Z(
        n5499) );
  HS65_LS_AOI212X2 U11230 ( .A(n710), .B(n679), .C(n676), .D(n711), .E(n5504), 
        .Z(n5501) );
  HS65_LS_NAND2X2 U11231 ( .A(n447), .B(n423), .Z(n3817) );
  HS65_LS_NOR4ABX2 U11232 ( .A(n7780), .B(n8865), .C(n8866), .D(n8867), .Z(
        n8864) );
  HS65_LS_MX41X4 U11233 ( .D0(n335), .S0(n356), .D1(n326), .S1(n353), .D2(n341), .S2(n332), .D3(n329), .S3(n349), .Z(n8866) );
  HS65_LS_NOR4ABX2 U11234 ( .A(n7763), .B(n8656), .C(n8657), .D(n8658), .Z(
        n8655) );
  HS65_LS_MX41X4 U11235 ( .D0(n370), .S0(n394), .D1(n377), .S1(n396), .D2(n403), .S2(n381), .D3(n378), .S3(n390), .Z(n8657) );
  HS65_LS_NAND4ABX3 U11236 ( .A(n8338), .B(n8339), .C(n8340), .D(n8341), .Z(
        n8055) );
  HS65_LS_NAND4ABX3 U11237 ( .A(n8367), .B(n8368), .C(n8369), .D(n8370), .Z(
        n8339) );
  HS65_LS_MX41X4 U11238 ( .D0(n318), .S0(n353), .D1(n358), .S1(n321), .D2(n323), .S2(n348), .D3(n357), .S3(n329), .Z(n8338) );
  HS65_LS_NOR4ABX2 U11239 ( .A(n8342), .B(n8343), .C(n8344), .D(n8345), .Z(
        n8341) );
  HS65_LS_NAND2X2 U11240 ( .A(n192), .B(n225), .Z(n3509) );
  HS65_LS_NAND2X2 U11241 ( .A(n327), .B(n349), .Z(n8066) );
  HS65_LS_NAND2X2 U11242 ( .A(n365), .B(n387), .Z(n8121) );
  HS65_LS_NAND2X2 U11243 ( .A(n598), .B(n611), .Z(n8690) );
  HS65_LS_NAND2X2 U11244 ( .A(n111), .B(n124), .Z(n8778) );
  HS65_LS_NAND4ABX3 U11245 ( .A(n3630), .B(n3631), .C(n3632), .D(n3633), .Z(
        n3249) );
  HS65_LS_NOR4ABX2 U11246 ( .A(n3634), .B(n3635), .C(n3636), .D(n3637), .Z(
        n3633) );
  HS65_LS_NAND3AX3 U11247 ( .A(n3642), .B(n3643), .C(n3644), .Z(n3631) );
  HS65_LS_NAND4ABX3 U11248 ( .A(n3646), .B(n3647), .C(n3648), .D(n3649), .Z(
        n3630) );
  HS65_LS_NAND4ABX3 U11249 ( .A(n2445), .B(n2446), .C(n2447), .D(n2448), .Z(
        n2358) );
  HS65_LS_NOR4ABX2 U11250 ( .A(n2449), .B(n2450), .C(n2451), .D(n2265), .Z(
        n2448) );
  HS65_LS_NOR3AX2 U11251 ( .A(n2452), .B(n2453), .C(n2454), .Z(n2447) );
  HS65_LS_NAND4ABX3 U11252 ( .A(n2460), .B(n2461), .C(n2462), .D(n2463), .Z(
        n2445) );
  HS65_LS_NAND4ABX3 U11253 ( .A(n1693), .B(n1694), .C(n1695), .D(n1696), .Z(
        n1606) );
  HS65_LS_NOR4ABX2 U11254 ( .A(n1697), .B(n1698), .C(n1699), .D(n1513), .Z(
        n1696) );
  HS65_LS_NOR3AX2 U11255 ( .A(n1700), .B(n1701), .C(n1702), .Z(n1695) );
  HS65_LS_NAND4ABX3 U11256 ( .A(n1708), .B(n1709), .C(n1710), .D(n1711), .Z(
        n1693) );
  HS65_LS_NAND4ABX3 U11257 ( .A(n1317), .B(n1318), .C(n1319), .D(n1320), .Z(
        n1230) );
  HS65_LS_NOR4ABX2 U11258 ( .A(n1321), .B(n1322), .C(n1323), .D(n1137), .Z(
        n1320) );
  HS65_LS_NOR3AX2 U11259 ( .A(n1324), .B(n1325), .C(n1326), .Z(n1319) );
  HS65_LS_NAND4ABX3 U11260 ( .A(n1332), .B(n1333), .C(n1334), .D(n1335), .Z(
        n1317) );
  HS65_LS_NAND4ABX3 U11261 ( .A(n2069), .B(n2070), .C(n2071), .D(n2072), .Z(
        n1982) );
  HS65_LS_NOR4ABX2 U11262 ( .A(n2073), .B(n2074), .C(n2075), .D(n1889), .Z(
        n2072) );
  HS65_LS_NOR3AX2 U11263 ( .A(n2076), .B(n2077), .C(n2078), .Z(n2071) );
  HS65_LS_NAND4ABX3 U11264 ( .A(n2084), .B(n2085), .C(n2086), .D(n2087), .Z(
        n2069) );
  HS65_LS_NAND4ABX3 U11265 ( .A(n3850), .B(n3851), .C(n3852), .D(n3853), .Z(
        n3378) );
  HS65_LS_NOR3AX2 U11266 ( .A(n3857), .B(n3858), .C(n3859), .Z(n3852) );
  HS65_LS_NOR4ABX2 U11267 ( .A(n3854), .B(n3855), .C(n3856), .D(n2857), .Z(
        n3853) );
  HS65_LS_NAND4ABX3 U11268 ( .A(n3865), .B(n3866), .C(n3867), .D(n3868), .Z(
        n3850) );
  HS65_LS_NAND3X2 U11269 ( .A(n8840), .B(n8841), .C(n8842), .Z(n8462) );
  HS65_LS_NOR4ABX2 U11270 ( .A(n8847), .B(n7742), .C(n7902), .D(n8848), .Z(
        n8841) );
  HS65_LS_NOR4ABX2 U11271 ( .A(n8849), .B(n7937), .C(n8850), .D(n8851), .Z(
        n8840) );
  HS65_LS_NOR4ABX2 U11272 ( .A(n7924), .B(n8843), .C(n8844), .D(n8845), .Z(
        n8842) );
  HS65_LS_NAND4ABX3 U11273 ( .A(n3491), .B(n3492), .C(n3493), .D(n3494), .Z(
        n3087) );
  HS65_LS_NOR3AX2 U11274 ( .A(n3499), .B(n3500), .C(n3501), .Z(n3493) );
  HS65_LS_NAND4ABX3 U11275 ( .A(n3503), .B(n3504), .C(n3505), .D(n3506), .Z(
        n3492) );
  HS65_LS_NOR4ABX2 U11276 ( .A(n3495), .B(n3496), .C(n3497), .D(n3498), .Z(
        n3494) );
  HS65_LS_NOR4ABX2 U11277 ( .A(n2343), .B(n2294), .C(n2278), .D(n2357), .Z(
        n2396) );
  HS65_LS_NOR4ABX2 U11278 ( .A(n1215), .B(n1166), .C(n1150), .D(n1229), .Z(
        n1268) );
  HS65_LS_NOR4ABX2 U11279 ( .A(n1967), .B(n1918), .C(n1902), .D(n1981), .Z(
        n2020) );
  HS65_LS_NOR4ABX2 U11280 ( .A(n1591), .B(n1542), .C(n1526), .D(n1605), .Z(
        n1644) );
  HS65_LS_NAND4ABX3 U11281 ( .A(n3733), .B(n3734), .C(n3735), .D(n3736), .Z(
        n3316) );
  HS65_LS_NAND4ABX3 U11282 ( .A(n3744), .B(n3745), .C(n3746), .D(n3747), .Z(
        n3734) );
  HS65_LS_NOR4ABX2 U11283 ( .A(n3737), .B(n3738), .C(n3739), .D(n2902), .Z(
        n3736) );
  HS65_LS_NOR3AX2 U11284 ( .A(n3740), .B(n3741), .C(n3742), .Z(n3735) );
  HS65_LS_NAND4ABX3 U11285 ( .A(n8271), .B(n8272), .C(n8273), .D(n8274), .Z(
        n8105) );
  HS65_LS_NOR4ABX2 U11286 ( .A(n8275), .B(n8276), .C(n8277), .D(n8278), .Z(
        n8274) );
  HS65_LS_OR4X4 U11287 ( .A(n8287), .B(n7756), .C(n8288), .D(n8289), .Z(n8271)
         );
  HS65_LS_NAND3AX3 U11288 ( .A(n8283), .B(n8284), .C(n8285), .Z(n8272) );
  HS65_LS_NOR4ABX2 U11289 ( .A(n3076), .B(n2867), .C(n2937), .D(n3086), .Z(
        n3424) );
  HS65_LS_NOR4ABX2 U11290 ( .A(n3305), .B(n2979), .C(n3140), .D(n3315), .Z(
        n3668) );
  HS65_LS_NOR4ABX2 U11291 ( .A(n3367), .B(n2997), .C(n3181), .D(n3377), .Z(
        n3785) );
  HS65_LS_NAND4ABX3 U11292 ( .A(n8704), .B(n8705), .C(n8706), .D(n8707), .Z(
        n8401) );
  HS65_LS_NOR4ABX2 U11293 ( .A(n7706), .B(n7647), .C(n7808), .D(n8708), .Z(
        n8707) );
  HS65_LS_NAND4ABX3 U11294 ( .A(n8715), .B(n7682), .C(n8716), .D(n7826), .Z(
        n8704) );
  HS65_LS_NOR4ABX2 U11295 ( .A(n8709), .B(n8710), .C(n7837), .D(n8711), .Z(
        n8706) );
  HS65_LS_NAND4ABX3 U11296 ( .A(n8792), .B(n8793), .C(n8794), .D(n8795), .Z(
        n8461) );
  HS65_LS_NOR4ABX2 U11297 ( .A(n7744), .B(n7675), .C(n7908), .D(n8796), .Z(
        n8795) );
  HS65_LS_NAND4ABX3 U11298 ( .A(n8803), .B(n7720), .C(n8804), .D(n7925), .Z(
        n8792) );
  HS65_LS_NOR4ABX2 U11299 ( .A(n8797), .B(n8798), .C(n7936), .D(n8799), .Z(
        n8794) );
  HS65_LS_NOR4ABX2 U11300 ( .A(n4105), .B(n4091), .C(n3997), .D(n4138), .Z(
        n4137) );
  HS65_LS_MX41X4 U11301 ( .D0(n148), .S0(n175), .D1(n170), .S1(n159), .D2(n165), .S2(n155), .D3(n154), .S3(n181), .Z(n4138) );
  HS65_LS_NAND2X2 U11302 ( .A(n375), .B(n390), .Z(n8023) );
  HS65_LS_NOR4ABX2 U11303 ( .A(n6915), .B(n6904), .C(n6925), .D(n6884), .Z(
        n7452) );
  HS65_LS_NOR4ABX2 U11304 ( .A(n5438), .B(n5427), .C(n5448), .D(n5407), .Z(
        n5919) );
  HS65_LS_NOR4ABX2 U11305 ( .A(n7030), .B(n7019), .C(n7040), .D(n6999), .Z(
        n7511) );
  HS65_LS_NOR4ABX2 U11306 ( .A(n5323), .B(n5312), .C(n5333), .D(n5292), .Z(
        n5860) );
  HS65_LS_NOR4ABX2 U11307 ( .A(n5207), .B(n5196), .C(n5217), .D(n5175), .Z(
        n5702) );
  HS65_LS_NOR4ABX2 U11308 ( .A(n6799), .B(n6788), .C(n6809), .D(n6767), .Z(
        n7294) );
  HS65_LS_NOR4ABX2 U11309 ( .A(n2147), .B(n2148), .C(n2149), .D(n2150), .Z(
        n2146) );
  HS65_LS_MX41X4 U11310 ( .D0(n787), .S0(n797), .D1(n799), .S1(n777), .D2(n772), .S2(n798), .D3(n804), .S3(n775), .Z(n2150) );
  HS65_LS_NOR4ABX2 U11311 ( .A(n1395), .B(n1396), .C(n1397), .D(n1398), .Z(
        n1394) );
  HS65_LS_MX41X4 U11312 ( .D0(n869), .S0(n879), .D1(n881), .S1(n859), .D2(n854), .S2(n880), .D3(n886), .S3(n857), .Z(n1398) );
  HS65_LS_NOR4ABX2 U11313 ( .A(n1771), .B(n1772), .C(n1773), .D(n1774), .Z(
        n1770) );
  HS65_LS_MX41X4 U11314 ( .D0(n828), .S0(n838), .D1(n840), .S1(n818), .D2(n813), .S2(n839), .D3(n845), .S3(n816), .Z(n1774) );
  HS65_LS_NOR4ABX2 U11315 ( .A(n2523), .B(n2524), .C(n2525), .D(n2526), .Z(
        n2522) );
  HS65_LS_MX41X4 U11316 ( .D0(n910), .S0(n920), .D1(n922), .S1(n900), .D2(n895), .S2(n921), .D3(n927), .S3(n898), .Z(n2526) );
  HS65_LS_NOR4ABX2 U11317 ( .A(n7636), .B(n7689), .C(n9014), .D(n7702), .Z(
        n9013) );
  HS65_LS_MX41X4 U11318 ( .D0(n619), .S0(n585), .D1(n614), .S1(n598), .D2(n623), .S2(n593), .D3(n594), .S3(n611), .Z(n9014) );
  HS65_LS_NOR4ABX2 U11319 ( .A(n7664), .B(n7727), .C(n9072), .D(n7740), .Z(
        n9071) );
  HS65_LS_MX41X4 U11320 ( .D0(n132), .S0(n98), .D1(n127), .S1(n111), .D2(n136), 
        .S2(n106), .D3(n107), .S3(n124), .Z(n9072) );
  HS65_LS_NAND2X2 U11321 ( .A(n76), .B(n56), .Z(n6850) );
  HS65_LS_NAND2X2 U11322 ( .A(n255), .B(n235), .Z(n5258) );
  HS65_LS_NAND2X2 U11323 ( .A(n474), .B(n454), .Z(n5373) );
  HS65_LS_NAND2X2 U11324 ( .A(n297), .B(n277), .Z(n6965) );
  HS65_LS_NAND2X2 U11325 ( .A(n528), .B(n506), .Z(n6732) );
  HS65_LS_NAND2X2 U11326 ( .A(n710), .B(n688), .Z(n5140) );
  HS65_LS_NOR4ABX2 U11327 ( .A(n5561), .B(n5562), .C(n5563), .D(n5564), .Z(
        n5560) );
  HS65_LS_MX41X4 U11328 ( .D0(n461), .S0(n486), .D1(n460), .S1(n483), .D2(n479), .S2(n455), .D3(n454), .S3(n471), .Z(n5563) );
  HS65_LS_NOR4ABX2 U11329 ( .A(n5540), .B(n5541), .C(n5542), .D(n5543), .Z(
        n5539) );
  HS65_LS_MX41X4 U11330 ( .D0(n242), .S0(n267), .D1(n241), .S1(n264), .D2(n260), .S2(n236), .D3(n235), .S3(n252), .Z(n5542) );
  HS65_LS_NOR4ABX2 U11331 ( .A(n7153), .B(n7154), .C(n7155), .D(n7156), .Z(
        n7152) );
  HS65_LS_MX41X4 U11332 ( .D0(n284), .S0(n309), .D1(n283), .S1(n306), .D2(n302), .S2(n278), .D3(n277), .S3(n294), .Z(n7155) );
  HS65_LS_NOR4ABX2 U11333 ( .A(n5684), .B(n5578), .C(n5793), .D(n5704), .Z(
        n5792) );
  HS65_LS_MX41X4 U11334 ( .D0(n679), .S0(n705), .D1(n686), .S1(n701), .D2(n693), .S2(n689), .D3(n688), .S3(n711), .Z(n5793) );
  HS65_LS_NOR4ABX2 U11335 ( .A(n5654), .B(n5513), .C(n5731), .D(n5674), .Z(
        n5730) );
  HS65_LS_MX41X4 U11336 ( .D0(n14), .S0(n41), .D1(n22), .S1(n37), .D2(n25), 
        .S2(n29), .D3(n24), .S3(n47), .Z(n5731) );
  HS65_LS_NOR4ABX2 U11337 ( .A(n7276), .B(n7170), .C(n7385), .D(n7296), .Z(
        n7384) );
  HS65_LS_MX41X4 U11338 ( .D0(n497), .S0(n523), .D1(n504), .S1(n519), .D2(n511), .S2(n507), .D3(n506), .S3(n529), .Z(n7385) );
  HS65_LS_NOR4ABX2 U11339 ( .A(n7132), .B(n7133), .C(n7134), .D(n7135), .Z(
        n7131) );
  HS65_LS_MX41X4 U11340 ( .D0(n63), .S0(n88), .D1(n62), .S1(n85), .D2(n81), 
        .S2(n57), .D3(n56), .S3(n73), .Z(n7134) );
  HS65_LS_NOR4ABX2 U11341 ( .A(n7246), .B(n7105), .C(n7323), .D(n7266), .Z(
        n7322) );
  HS65_LS_MX41X4 U11342 ( .D0(n540), .S0(n567), .D1(n548), .S1(n563), .D2(n551), .S2(n555), .D3(n550), .S3(n573), .Z(n7323) );
  HS65_LS_NAND4ABX3 U11343 ( .A(n9032), .B(n9033), .C(n9034), .D(n9035), .Z(
        n7701) );
  HS65_LS_AOI222X2 U11344 ( .A(n591), .B(n623), .C(n594), .D(n613), .E(n598), 
        .F(n624), .Z(n9034) );
  HS65_LS_NAND4ABX3 U11345 ( .A(n588), .B(n8760), .C(n8696), .D(n8407), .Z(
        n9033) );
  HS65_LS_NOR4ABX2 U11346 ( .A(n8731), .B(n8724), .C(n8739), .D(n8708), .Z(
        n9035) );
  HS65_LS_NAND4ABX3 U11347 ( .A(n9090), .B(n9091), .C(n9092), .D(n9093), .Z(
        n7739) );
  HS65_LS_AOI222X2 U11348 ( .A(n104), .B(n136), .C(n107), .D(n126), .E(n111), 
        .F(n137), .Z(n9092) );
  HS65_LS_NAND4ABX3 U11349 ( .A(n101), .B(n8848), .C(n8784), .D(n8467), .Z(
        n9091) );
  HS65_LS_NOR4ABX2 U11350 ( .A(n8819), .B(n8812), .C(n8827), .D(n8796), .Z(
        n9093) );
  HS65_LS_IVX2 U11351 ( .A(n3427), .Z(n196) );
  HS65_LS_NOR3AX2 U11352 ( .A(n3428), .B(n3429), .C(n3430), .Z(n3427) );
  HS65_LS_NOR4ABX2 U11353 ( .A(n6643), .B(n6668), .C(n6676), .D(n6688), .Z(
        n7264) );
  HS65_LS_NOR4ABX2 U11354 ( .A(n5050), .B(n5075), .C(n5083), .D(n5095), .Z(
        n5672) );
  HS65_LS_NOR4ABX2 U11355 ( .A(n3657), .B(n3606), .C(n3618), .D(n3647), .Z(
        n4102) );
  HS65_LS_IVX2 U11356 ( .A(n2794), .Z(n51) );
  HS65_LS_IVX2 U11357 ( .A(n2907), .Z(n142) );
  HS65_LS_NOR4ABX2 U11358 ( .A(n8579), .B(n8580), .C(n8581), .D(n8582), .Z(
        n8578) );
  HS65_LS_NAND2X2 U11359 ( .A(n633), .B(n663), .Z(n3347) );
  HS65_LS_NAND3X2 U11360 ( .A(n8896), .B(n8897), .C(n8898), .Z(n8867) );
  HS65_LS_NOR4X4 U11361 ( .A(n8526), .B(n8382), .C(n8367), .D(n8356), .Z(n8897) );
  HS65_LS_NOR4ABX2 U11362 ( .A(n8602), .B(n8066), .C(n8899), .D(n8900), .Z(
        n8898) );
  HS65_LS_NOR4ABX2 U11363 ( .A(n8552), .B(n7966), .C(n8564), .D(n8537), .Z(
        n8896) );
  HS65_LS_NAND2X2 U11364 ( .A(n358), .B(n318), .Z(n8529) );
  HS65_LS_NOR4ABX2 U11365 ( .A(n6647), .B(n6648), .C(n6649), .D(n6650), .Z(
        n6641) );
  HS65_LS_NOR4ABX2 U11366 ( .A(n5054), .B(n5055), .C(n5056), .D(n5057), .Z(
        n5048) );
  HS65_LS_NOR4ABX2 U11367 ( .A(n6707), .B(n6708), .C(n6709), .D(n6710), .Z(
        n6275) );
  HS65_LS_NAND3AX3 U11368 ( .A(n6711), .B(n6712), .C(n6713), .Z(n6710) );
  HS65_LS_NAND4ABX3 U11369 ( .A(n6714), .B(n6715), .C(n6716), .D(n6717), .Z(
        n6709) );
  HS65_LS_AOI212X2 U11370 ( .A(n540), .B(n6718), .C(n569), .D(n6719), .E(n6720), .Z(n6708) );
  HS65_LS_NOR4ABX2 U11371 ( .A(n5114), .B(n5115), .C(n5116), .D(n5117), .Z(
        n4682) );
  HS65_LS_NAND3AX3 U11372 ( .A(n5118), .B(n5119), .C(n5120), .Z(n5117) );
  HS65_LS_NAND4ABX3 U11373 ( .A(n5121), .B(n5122), .C(n5123), .D(n5124), .Z(
        n5116) );
  HS65_LS_AOI212X2 U11374 ( .A(n14), .B(n5125), .C(n43), .D(n5126), .E(n5127), 
        .Z(n5115) );
  HS65_LS_NAND2X2 U11375 ( .A(n159), .B(n171), .Z(n3062) );
  HS65_LS_NAND3X2 U11376 ( .A(n8956), .B(n8957), .C(n8958), .Z(n8658) );
  HS65_LS_NOR4X4 U11377 ( .A(n8221), .B(n8088), .C(n8125), .D(n8114), .Z(n8957) );
  HS65_LS_NOR4ABX2 U11378 ( .A(n8248), .B(n7864), .C(n8260), .D(n8310), .Z(
        n8956) );
  HS65_LS_NOR4ABX2 U11379 ( .A(n8298), .B(n8023), .C(n8959), .D(n8960), .Z(
        n8958) );
  HS65_LS_NOR4ABX2 U11380 ( .A(n3534), .B(n2953), .C(n3094), .D(n3464), .Z(
        n4204) );
  HS65_LS_IVX2 U11381 ( .A(n2745), .Z(n630) );
  HS65_LS_NOR4ABX2 U11382 ( .A(n8115), .B(n8116), .C(n8117), .D(n8118), .Z(
        n8109) );
  HS65_LS_NAND2X2 U11383 ( .A(n144), .B(n179), .Z(n2930) );
  HS65_LS_NOR4ABX2 U11384 ( .A(n8353), .B(n8354), .C(n8355), .D(n8356), .Z(
        n8352) );
  HS65_LS_NOR4ABX2 U11385 ( .A(n6941), .B(n6942), .C(n6943), .D(n6944), .Z(
        n6514) );
  HS65_LS_NAND3AX3 U11386 ( .A(n6945), .B(n6946), .C(n6947), .Z(n6943) );
  HS65_LS_NOR4ABX2 U11387 ( .A(n6953), .B(n6954), .C(n6955), .D(n6956), .Z(
        n6941) );
  HS65_LS_MX41X4 U11388 ( .D0(n66), .S0(n91), .D1(n76), .S1(n59), .D2(n81), 
        .S2(n65), .D3(n86), .S3(n60), .Z(n6944) );
  HS65_LS_NOR4ABX2 U11389 ( .A(n7056), .B(n7057), .C(n7058), .D(n7059), .Z(
        n6568) );
  HS65_LS_NAND3AX3 U11390 ( .A(n7060), .B(n7061), .C(n7062), .Z(n7058) );
  HS65_LS_NOR4ABX2 U11391 ( .A(n7068), .B(n7069), .C(n7070), .D(n7071), .Z(
        n7056) );
  HS65_LS_MX41X4 U11392 ( .D0(n287), .S0(n312), .D1(n297), .S1(n280), .D2(n302), .S2(n286), .D3(n307), .S3(n281), .Z(n7059) );
  HS65_LS_NOR4ABX2 U11393 ( .A(n5464), .B(n5465), .C(n5466), .D(n5467), .Z(
        n4975) );
  HS65_LS_NAND3AX3 U11394 ( .A(n5468), .B(n5469), .C(n5470), .Z(n5466) );
  HS65_LS_NOR4ABX2 U11395 ( .A(n5476), .B(n5477), .C(n5478), .D(n5479), .Z(
        n5464) );
  HS65_LS_MX41X4 U11396 ( .D0(n464), .S0(n489), .D1(n474), .S1(n457), .D2(n479), .S2(n463), .D3(n484), .S3(n458), .Z(n5467) );
  HS65_LS_NOR4ABX2 U11397 ( .A(n5349), .B(n5350), .C(n5351), .D(n5352), .Z(
        n4921) );
  HS65_LS_NAND3AX3 U11398 ( .A(n5353), .B(n5354), .C(n5355), .Z(n5351) );
  HS65_LS_NOR4ABX2 U11399 ( .A(n5361), .B(n5362), .C(n5363), .D(n5364), .Z(
        n5349) );
  HS65_LS_MX41X4 U11400 ( .D0(n245), .S0(n270), .D1(n255), .S1(n238), .D2(n260), .S2(n244), .D3(n265), .S3(n239), .Z(n5352) );
  HS65_LS_NOR4ABX2 U11401 ( .A(n5234), .B(n5235), .C(n5236), .D(n5237), .Z(
        n4845) );
  HS65_LS_NAND3AX3 U11402 ( .A(n5238), .B(n5239), .C(n5240), .Z(n5236) );
  HS65_LS_NOR4ABX2 U11403 ( .A(n5246), .B(n5247), .C(n5248), .D(n5249), .Z(
        n5234) );
  HS65_LS_MX41X4 U11404 ( .D0(n680), .S0(n706), .D1(n710), .S1(n684), .D2(n693), .S2(n682), .D3(n699), .S3(n683), .Z(n5237) );
  HS65_LS_NOR4ABX2 U11405 ( .A(n6826), .B(n6827), .C(n6828), .D(n6829), .Z(
        n6438) );
  HS65_LS_NAND3AX3 U11406 ( .A(n6830), .B(n6831), .C(n6832), .Z(n6828) );
  HS65_LS_NOR4ABX2 U11407 ( .A(n6838), .B(n6839), .C(n6840), .D(n6841), .Z(
        n6826) );
  HS65_LS_MX41X4 U11408 ( .D0(n498), .S0(n524), .D1(n528), .S1(n502), .D2(n511), .S2(n500), .D3(n517), .S3(n501), .Z(n6829) );
  HS65_LS_NOR4ABX2 U11409 ( .A(n8610), .B(n8611), .C(n8612), .D(n8613), .Z(
        n8347) );
  HS65_LS_MX41X4 U11410 ( .D0(n334), .S0(n354), .D1(n323), .S1(n347), .D2(n341), .S2(n336), .D3(n324), .S3(n350), .Z(n8613) );
  HS65_LS_NAND4ABX3 U11411 ( .A(n8614), .B(n8615), .C(n8616), .D(n8617), .Z(
        n8612) );
  HS65_LS_NOR4ABX2 U11412 ( .A(n8622), .B(n8623), .C(n8624), .D(n8625), .Z(
        n8610) );
  HS65_LS_NOR4ABX2 U11413 ( .A(n3588), .B(n3589), .C(n3590), .D(n3591), .Z(
        n3029) );
  HS65_LS_NAND4ABX3 U11414 ( .A(n3592), .B(n3593), .C(n3594), .D(n3595), .Z(
        n3591) );
  HS65_LS_AOI212X2 U11415 ( .A(n180), .B(n3596), .C(n169), .D(n3597), .E(n3598), .Z(n3589) );
  HS65_LS_MX41X4 U11416 ( .D0(n155), .S0(n182), .D1(n160), .S1(n166), .D2(n172), .S2(n147), .D3(n177), .S3(n153), .Z(n3590) );
  HS65_LS_NOR4ABX2 U11417 ( .A(n1717), .B(n1673), .C(n1689), .D(n1708), .Z(
        n1823) );
  HS65_LS_NOR4ABX2 U11418 ( .A(n2469), .B(n2425), .C(n2441), .D(n2460), .Z(
        n2575) );
  HS65_LS_NAND2X2 U11419 ( .A(n106), .B(n126), .Z(n8837) );
  HS65_LS_NAND2X2 U11420 ( .A(n593), .B(n613), .Z(n8749) );
  HS65_LS_NAND2X2 U11421 ( .A(n36), .B(n26), .Z(n4730) );
  HS65_LS_NAND2X2 U11422 ( .A(n562), .B(n552), .Z(n6323) );
  HS65_LS_NOR4ABX2 U11423 ( .A(n1341), .B(n1297), .C(n1313), .D(n1332), .Z(
        n1447) );
  HS65_LS_NOR4ABX2 U11424 ( .A(n2093), .B(n2049), .C(n2065), .D(n2084), .Z(
        n2199) );
  HS65_LS_NOR4ABX2 U11425 ( .A(n2367), .B(n2368), .C(n2369), .D(n2370), .Z(
        n2361) );
  HS65_LS_NOR4ABX2 U11426 ( .A(n1615), .B(n1616), .C(n1617), .D(n1618), .Z(
        n1609) );
  HS65_LS_NAND2X2 U11427 ( .A(n481), .B(n456), .Z(n4998) );
  HS65_LS_NAND2X2 U11428 ( .A(n262), .B(n237), .Z(n4944) );
  HS65_LS_NAND2X2 U11429 ( .A(n304), .B(n279), .Z(n6591) );
  HS65_LS_NAND2X2 U11430 ( .A(n83), .B(n58), .Z(n6537) );
  HS65_LS_NAND2X2 U11431 ( .A(n700), .B(n690), .Z(n4870) );
  HS65_LS_NAND2X2 U11432 ( .A(n518), .B(n508), .Z(n6463) );
  HS65_LS_NOR4ABX2 U11433 ( .A(n3874), .B(n3830), .C(n3846), .D(n3865), .Z(
        n4310) );
  HS65_LS_NOR4ABX2 U11434 ( .A(n4268), .B(n3338), .C(n3763), .D(n3681), .Z(
        n4267) );
  HS65_LS_OAI21X2 U11435 ( .A(n646), .B(n647), .C(n661), .Z(n4268) );
  HS65_LS_NOR4ABX2 U11436 ( .A(n3662), .B(n3616), .C(n3605), .D(n3641), .Z(
        n4132) );
  HS65_LS_NAND2X2 U11437 ( .A(n903), .B(n922), .Z(n2320) );
  HS65_LS_NAND2X2 U11438 ( .A(n821), .B(n840), .Z(n1568) );
  HS65_LS_NOR4ABX2 U11439 ( .A(n3757), .B(n3713), .C(n3729), .D(n3748), .Z(
        n4251) );
  HS65_LS_NAND4ABX3 U11440 ( .A(n6493), .B(n6494), .C(n6495), .D(n6496), .Z(
        n6190) );
  HS65_LS_NOR3X1 U11441 ( .A(n6497), .B(n6498), .C(n6499), .Z(n6496) );
  HS65_LS_AOI222X2 U11442 ( .A(n63), .B(n85), .C(n66), .D(n89), .E(n77), .F(
        n64), .Z(n6495) );
  HS65_LS_NAND3X2 U11443 ( .A(n6500), .B(n6501), .C(n6502), .Z(n6494) );
  HS65_LS_NAND4ABX3 U11444 ( .A(n6547), .B(n6548), .C(n6549), .D(n6550), .Z(
        n6202) );
  HS65_LS_NOR3X1 U11445 ( .A(n6551), .B(n6552), .C(n6553), .Z(n6550) );
  HS65_LS_AOI222X2 U11446 ( .A(n284), .B(n306), .C(n287), .D(n310), .E(n298), 
        .F(n285), .Z(n6549) );
  HS65_LS_NAND3X2 U11447 ( .A(n6554), .B(n6555), .C(n6556), .Z(n6548) );
  HS65_LS_NAND4ABX3 U11448 ( .A(n4900), .B(n4901), .C(n4902), .D(n4903), .Z(
        n4597) );
  HS65_LS_NOR3X1 U11449 ( .A(n4904), .B(n4905), .C(n4906), .Z(n4903) );
  HS65_LS_AOI222X2 U11450 ( .A(n242), .B(n264), .C(n245), .D(n268), .E(n256), 
        .F(n243), .Z(n4902) );
  HS65_LS_NAND3X2 U11451 ( .A(n4907), .B(n4908), .C(n4909), .Z(n4901) );
  HS65_LS_NAND4ABX3 U11452 ( .A(n4954), .B(n4955), .C(n4956), .D(n4957), .Z(
        n4609) );
  HS65_LS_NOR3X1 U11453 ( .A(n4958), .B(n4959), .C(n4960), .Z(n4957) );
  HS65_LS_AOI222X2 U11454 ( .A(n461), .B(n483), .C(n464), .D(n487), .E(n475), 
        .F(n462), .Z(n4956) );
  HS65_LS_NAND3X2 U11455 ( .A(n4961), .B(n4962), .C(n4963), .Z(n4955) );
  HS65_LS_NAND4ABX3 U11456 ( .A(n4823), .B(n4824), .C(n4825), .D(n4826), .Z(
        n4539) );
  HS65_LS_NOR3X1 U11457 ( .A(n4827), .B(n4828), .C(n4829), .Z(n4826) );
  HS65_LS_AOI222X2 U11458 ( .A(n679), .B(n701), .C(n680), .D(n704), .E(n709), 
        .F(n681), .Z(n4825) );
  HS65_LS_NAND3X2 U11459 ( .A(n4830), .B(n4831), .C(n4832), .Z(n4824) );
  HS65_LS_NAND4ABX3 U11460 ( .A(n6416), .B(n6417), .C(n6418), .D(n6419), .Z(
        n6132) );
  HS65_LS_NOR3X1 U11461 ( .A(n6420), .B(n6421), .C(n6422), .Z(n6419) );
  HS65_LS_AOI222X2 U11462 ( .A(n497), .B(n519), .C(n498), .D(n522), .E(n527), 
        .F(n499), .Z(n6418) );
  HS65_LS_NAND3X2 U11463 ( .A(n6423), .B(n6424), .C(n6425), .Z(n6417) );
  HS65_LS_NAND4ABX3 U11464 ( .A(n4683), .B(n4684), .C(n4685), .D(n4686), .Z(
        n4483) );
  HS65_LS_NOR3X1 U11465 ( .A(n4687), .B(n4688), .C(n4689), .Z(n4686) );
  HS65_LS_AOI222X2 U11466 ( .A(n14), .B(n37), .C(n40), .D(n15), .E(n45), .F(
        n16), .Z(n4685) );
  HS65_LS_NAND3X2 U11467 ( .A(n4690), .B(n4691), .C(n4692), .Z(n4684) );
  HS65_LS_NAND4ABX3 U11468 ( .A(n6276), .B(n6277), .C(n6278), .D(n6279), .Z(
        n6076) );
  HS65_LS_NOR3X1 U11469 ( .A(n6280), .B(n6281), .C(n6282), .Z(n6279) );
  HS65_LS_AOI222X2 U11470 ( .A(n540), .B(n563), .C(n566), .D(n541), .E(n571), 
        .F(n542), .Z(n6278) );
  HS65_LS_NAND3X2 U11471 ( .A(n6283), .B(n6284), .C(n6285), .Z(n6277) );
  HS65_LS_NAND2X2 U11472 ( .A(n862), .B(n881), .Z(n1192) );
  HS65_LS_NAND2X2 U11473 ( .A(n780), .B(n799), .Z(n1944) );
  HS65_LS_NOR4ABX2 U11474 ( .A(n6928), .B(n6929), .C(n6930), .D(n6931), .Z(
        n6492) );
  HS65_LS_NAND3AX3 U11475 ( .A(n6932), .B(n6933), .C(n6934), .Z(n6931) );
  HS65_LS_NAND4ABX3 U11476 ( .A(n6935), .B(n6936), .C(n6937), .D(n6938), .Z(
        n6930) );
  HS65_LS_AOI212X2 U11477 ( .A(n63), .B(n6939), .C(n87), .D(n6940), .E(n6067), 
        .Z(n6929) );
  HS65_LS_NOR4ABX2 U11478 ( .A(n5336), .B(n5337), .C(n5338), .D(n5339), .Z(
        n4899) );
  HS65_LS_NAND3AX3 U11479 ( .A(n5340), .B(n5341), .C(n5342), .Z(n5339) );
  HS65_LS_NAND4ABX3 U11480 ( .A(n5343), .B(n5344), .C(n5345), .D(n5346), .Z(
        n5338) );
  HS65_LS_AOI212X2 U11481 ( .A(n242), .B(n5347), .C(n266), .D(n5348), .E(n4474), .Z(n5337) );
  HS65_LS_NOR4ABX2 U11482 ( .A(n5451), .B(n5452), .C(n5453), .D(n5454), .Z(
        n4953) );
  HS65_LS_NAND3AX3 U11483 ( .A(n5455), .B(n5456), .C(n5457), .Z(n5454) );
  HS65_LS_NAND4ABX3 U11484 ( .A(n5458), .B(n5459), .C(n5460), .D(n5461), .Z(
        n5453) );
  HS65_LS_AOI212X2 U11485 ( .A(n461), .B(n5462), .C(n485), .D(n5463), .E(n4520), .Z(n5452) );
  HS65_LS_NOR4ABX2 U11486 ( .A(n7043), .B(n7044), .C(n7045), .D(n7046), .Z(
        n6546) );
  HS65_LS_NAND3AX3 U11487 ( .A(n7047), .B(n7048), .C(n7049), .Z(n7046) );
  HS65_LS_NAND4ABX3 U11488 ( .A(n7050), .B(n7051), .C(n7052), .D(n7053), .Z(
        n7045) );
  HS65_LS_AOI212X2 U11489 ( .A(n284), .B(n7054), .C(n308), .D(n7055), .E(n6113), .Z(n7044) );
  HS65_LS_NOR4ABX2 U11490 ( .A(n6812), .B(n6813), .C(n6814), .D(n6815), .Z(
        n6415) );
  HS65_LS_NAND3AX3 U11491 ( .A(n6816), .B(n6817), .C(n6818), .Z(n6815) );
  HS65_LS_NAND4ABX3 U11492 ( .A(n6819), .B(n6820), .C(n6821), .D(n6822), .Z(
        n6814) );
  HS65_LS_AOI212X2 U11493 ( .A(n497), .B(n6823), .C(n525), .D(n6824), .E(n6825), .Z(n6813) );
  HS65_LS_NOR4ABX2 U11494 ( .A(n5220), .B(n5221), .C(n5222), .D(n5223), .Z(
        n4822) );
  HS65_LS_NAND3AX3 U11495 ( .A(n5224), .B(n5225), .C(n5226), .Z(n5223) );
  HS65_LS_NAND4ABX3 U11496 ( .A(n5227), .B(n5228), .C(n5229), .D(n5230), .Z(
        n5222) );
  HS65_LS_AOI212X2 U11497 ( .A(n679), .B(n5231), .C(n707), .D(n5232), .E(n5233), .Z(n5221) );
  HS65_LS_NAND2X2 U11498 ( .A(n145), .B(n167), .Z(n3562) );
  HS65_LS_OAI21X2 U11499 ( .A(n17), .B(n4693), .C(n47), .Z(n4692) );
  HS65_LS_OAI21X2 U11500 ( .A(n543), .B(n6286), .C(n573), .Z(n6285) );
  HS65_LS_NAND2X2 U11501 ( .A(n341), .B(n318), .Z(n8574) );
  HS65_LS_OAI21X2 U11502 ( .A(n65), .B(n6503), .C(n73), .Z(n6502) );
  HS65_LS_OAI21X2 U11503 ( .A(n286), .B(n6557), .C(n294), .Z(n6556) );
  HS65_LS_OAI21X2 U11504 ( .A(n244), .B(n4910), .C(n252), .Z(n4909) );
  HS65_LS_OAI21X2 U11505 ( .A(n463), .B(n4964), .C(n471), .Z(n4963) );
  HS65_LS_OAI21X2 U11506 ( .A(n682), .B(n4833), .C(n711), .Z(n4832) );
  HS65_LS_OAI21X2 U11507 ( .A(n500), .B(n6426), .C(n529), .Z(n6425) );
  HS65_LS_NOR4ABX2 U11508 ( .A(n8829), .B(n8830), .C(n8831), .D(n8832), .Z(
        n8451) );
  HS65_LS_NAND3AX3 U11509 ( .A(n8833), .B(n7918), .C(n8834), .Z(n8832) );
  HS65_LS_AOI212X2 U11510 ( .A(n98), .B(n8838), .C(n133), .D(n8839), .E(n7888), 
        .Z(n8830) );
  HS65_LS_NAND4ABX3 U11511 ( .A(n8835), .B(n8836), .C(n8837), .D(n7904), .Z(
        n8831) );
  HS65_LS_NOR4ABX2 U11512 ( .A(n8741), .B(n8742), .C(n8743), .D(n8744), .Z(
        n8391) );
  HS65_LS_NAND3AX3 U11513 ( .A(n8745), .B(n7819), .C(n8746), .Z(n8744) );
  HS65_LS_AOI212X2 U11514 ( .A(n585), .B(n8750), .C(n620), .D(n8751), .E(n7849), .Z(n8742) );
  HS65_LS_NAND4ABX3 U11515 ( .A(n8747), .B(n8748), .C(n8749), .D(n7804), .Z(
        n8743) );
  HS65_LS_NAND3X2 U11516 ( .A(n8752), .B(n8753), .C(n8754), .Z(n8402) );
  HS65_LS_NOR4ABX2 U11517 ( .A(n8759), .B(n7704), .C(n7802), .D(n8760), .Z(
        n8753) );
  HS65_LS_NOR4ABX2 U11518 ( .A(n8761), .B(n7838), .C(n8762), .D(n8763), .Z(
        n8752) );
  HS65_LS_NOR4ABX2 U11519 ( .A(n7825), .B(n8755), .C(n8756), .D(n8757), .Z(
        n8754) );
  HS65_LS_NOR4ABX2 U11520 ( .A(n6885), .B(n6886), .C(n6887), .D(n6888), .Z(
        n6879) );
  HS65_LS_NOR4ABX2 U11521 ( .A(n5293), .B(n5294), .C(n5295), .D(n5296), .Z(
        n5287) );
  HS65_LS_NOR4ABX2 U11522 ( .A(n5408), .B(n5409), .C(n5410), .D(n5411), .Z(
        n5402) );
  HS65_LS_NOR4ABX2 U11523 ( .A(n7000), .B(n7001), .C(n7002), .D(n7003), .Z(
        n6994) );
  HS65_LS_NOR4ABX2 U11524 ( .A(n5176), .B(n5177), .C(n5178), .D(n5179), .Z(
        n5170) );
  HS65_LS_NOR4ABX2 U11525 ( .A(n6768), .B(n6769), .C(n6770), .D(n6771), .Z(
        n6762) );
  HS65_LS_NOR4ABX2 U11526 ( .A(n3325), .B(n3326), .C(n3327), .D(n3328), .Z(
        n3319) );
  HS65_LS_NOR3AX2 U11527 ( .A(n7948), .B(n8055), .C(n8337), .Z(n8321) );
  HS65_LS_NAND2X2 U11528 ( .A(n391), .B(n375), .Z(n8284) );
  HS65_LS_NAND2X2 U11529 ( .A(n149), .B(n171), .Z(n3649) );
  HS65_LS_NOR4ABX2 U11530 ( .A(n5098), .B(n5099), .C(n5100), .D(n5101), .Z(
        n4705) );
  HS65_LS_NAND3AX3 U11531 ( .A(n5102), .B(n5103), .C(n5104), .Z(n5100) );
  HS65_LS_MX41X4 U11532 ( .D0(n42), .S0(n15), .D1(n46), .S1(n20), .D2(n17), 
        .S2(n29), .D3(n18), .S3(n35), .Z(n5101) );
  HS65_LS_NOR4ABX2 U11533 ( .A(n5110), .B(n5111), .C(n5112), .D(n5113), .Z(
        n5098) );
  HS65_LS_NOR4ABX2 U11534 ( .A(n6691), .B(n6692), .C(n6693), .D(n6694), .Z(
        n6298) );
  HS65_LS_NAND3AX3 U11535 ( .A(n6695), .B(n6696), .C(n6697), .Z(n6693) );
  HS65_LS_MX41X4 U11536 ( .D0(n568), .S0(n541), .D1(n572), .S1(n546), .D2(n543), .S2(n555), .D3(n544), .S3(n561), .Z(n6694) );
  HS65_LS_NOR4ABX2 U11537 ( .A(n6703), .B(n6704), .C(n6705), .D(n6706), .Z(
        n6691) );
  HS65_LS_NOR4ABX2 U11538 ( .A(n8279), .B(n8280), .C(n8281), .D(n8282), .Z(
        n8273) );
  HS65_LS_NAND2X2 U11539 ( .A(n172), .B(n153), .Z(n3624) );
  HS65_LS_NAND2X2 U11540 ( .A(n396), .B(n369), .Z(n8223) );
  HS65_LS_NAND4ABX3 U11541 ( .A(n4099), .B(n4100), .C(n4101), .D(n4102), .Z(
        n3923) );
  HS65_LS_NAND4ABX3 U11542 ( .A(n3287), .B(n3038), .C(n3272), .D(n3255), .Z(
        n4100) );
  HS65_LS_AOI222X2 U11543 ( .A(n143), .B(n165), .C(n154), .D(n172), .E(n166), 
        .F(n159), .Z(n4101) );
  HS65_LS_NAND4ABX3 U11544 ( .A(n3580), .B(n3592), .C(n4104), .D(n3562), .Z(
        n4099) );
  HS65_LS_NAND2X2 U11545 ( .A(n394), .B(n378), .Z(n8135) );
  HS65_LS_NAND4ABX3 U11546 ( .A(n1444), .B(n1445), .C(n1446), .D(n1447), .Z(
        n1387) );
  HS65_LS_AOI222X2 U11547 ( .A(n854), .B(n882), .C(n866), .D(n886), .E(n868), 
        .F(n881), .Z(n1446) );
  HS65_LS_NAND4ABX3 U11548 ( .A(n1260), .B(n1226), .C(n1183), .D(n1239), .Z(
        n1445) );
  HS65_LS_NAND4ABX3 U11549 ( .A(n1379), .B(n1367), .C(n1448), .D(n1284), .Z(
        n1444) );
  HS65_LS_NAND4ABX3 U11550 ( .A(n2196), .B(n2197), .C(n2198), .D(n2199), .Z(
        n2139) );
  HS65_LS_AOI222X2 U11551 ( .A(n772), .B(n800), .C(n784), .D(n804), .E(n786), 
        .F(n799), .Z(n2198) );
  HS65_LS_NAND4ABX3 U11552 ( .A(n2012), .B(n1978), .C(n1935), .D(n1991), .Z(
        n2197) );
  HS65_LS_NAND4ABX3 U11553 ( .A(n2131), .B(n2119), .C(n2200), .D(n2036), .Z(
        n2196) );
  HS65_LS_NAND4ABX3 U11554 ( .A(n1820), .B(n1821), .C(n1822), .D(n1823), .Z(
        n1763) );
  HS65_LS_AOI222X2 U11555 ( .A(n813), .B(n841), .C(n825), .D(n845), .E(n827), 
        .F(n840), .Z(n1822) );
  HS65_LS_NAND4ABX3 U11556 ( .A(n1755), .B(n1743), .C(n1824), .D(n1660), .Z(
        n1820) );
  HS65_LS_NAND4ABX3 U11557 ( .A(n1636), .B(n1602), .C(n1559), .D(n1615), .Z(
        n1821) );
  HS65_LS_NAND4ABX3 U11558 ( .A(n2572), .B(n2573), .C(n2574), .D(n2575), .Z(
        n2515) );
  HS65_LS_AOI222X2 U11559 ( .A(n895), .B(n923), .C(n907), .D(n927), .E(n909), 
        .F(n922), .Z(n2574) );
  HS65_LS_NAND4ABX3 U11560 ( .A(n2507), .B(n2495), .C(n2576), .D(n2412), .Z(
        n2572) );
  HS65_LS_NAND4ABX3 U11561 ( .A(n2388), .B(n2354), .C(n2311), .D(n2367), .Z(
        n2573) );
  HS65_LS_NAND2X2 U11562 ( .A(n175), .B(n152), .Z(n3607) );
  HS65_LS_NOR4ABX2 U11563 ( .A(n1621), .B(n1691), .C(n1716), .D(n1709), .Z(
        n1839) );
  HS65_LS_NOR4ABX2 U11564 ( .A(n2373), .B(n2443), .C(n2468), .D(n2461), .Z(
        n2591) );
  HS65_LS_NAND2X2 U11565 ( .A(n83), .B(n63), .Z(n6950) );
  HS65_LS_NAND2X2 U11566 ( .A(n481), .B(n461), .Z(n5473) );
  HS65_LS_NAND2X2 U11567 ( .A(n304), .B(n284), .Z(n7065) );
  HS65_LS_NAND2X2 U11568 ( .A(n262), .B(n242), .Z(n5358) );
  HS65_LS_NAND2X2 U11569 ( .A(n700), .B(n679), .Z(n5243) );
  HS65_LS_NAND2X2 U11570 ( .A(n518), .B(n497), .Z(n6835) );
  HS65_LS_OAI21X2 U11571 ( .A(n24), .B(n4693), .C(n42), .Z(n5491) );
  HS65_LS_OAI21X2 U11572 ( .A(n550), .B(n6286), .C(n568), .Z(n7083) );
  HS65_LS_OAI21X2 U11573 ( .A(n454), .B(n4964), .C(n489), .Z(n5570) );
  HS65_LS_OAI21X2 U11574 ( .A(n277), .B(n6557), .C(n312), .Z(n7162) );
  HS65_LS_OAI21X2 U11575 ( .A(n56), .B(n6503), .C(n91), .Z(n7141) );
  HS65_LS_OAI21X2 U11576 ( .A(n235), .B(n4910), .C(n270), .Z(n5549) );
  HS65_LS_NAND2X2 U11577 ( .A(n919), .B(n894), .Z(n2367) );
  HS65_LS_NAND2X2 U11578 ( .A(n837), .B(n812), .Z(n1615) );
  HS65_LS_NAND2X2 U11579 ( .A(n167), .B(n155), .Z(n3061) );
  HS65_LS_NAND2X2 U11580 ( .A(n878), .B(n853), .Z(n1239) );
  HS65_LS_NOR4ABX2 U11581 ( .A(n3638), .B(n3639), .C(n3640), .D(n3641), .Z(
        n3632) );
  HS65_LS_NAND2X2 U11582 ( .A(n399), .B(n377), .Z(n8008) );
  HS65_LS_NAND2X2 U11583 ( .A(n358), .B(n327), .Z(n8528) );
  HS65_LS_NAND2X2 U11584 ( .A(n796), .B(n771), .Z(n1991) );
  HS65_LS_NAND2X2 U11585 ( .A(n318), .B(n347), .Z(n8363) );
  HS65_LS_NAND2X2 U11586 ( .A(n147), .B(n180), .Z(n3255) );
  HS65_LS_NAND2X2 U11587 ( .A(n647), .B(n656), .Z(n3325) );
  HS65_LS_NAND2X2 U11588 ( .A(n86), .B(n63), .Z(n6500) );
  HS65_LS_NAND2X2 U11589 ( .A(n307), .B(n284), .Z(n6554) );
  HS65_LS_NAND2X2 U11590 ( .A(n265), .B(n242), .Z(n4907) );
  HS65_LS_NAND2X2 U11591 ( .A(n484), .B(n461), .Z(n4961) );
  HS65_LS_NAND2X2 U11592 ( .A(n699), .B(n679), .Z(n4830) );
  HS65_LS_NAND2X2 U11593 ( .A(n517), .B(n497), .Z(n6423) );
  HS65_LS_NAND2X2 U11594 ( .A(n145), .B(n169), .Z(n3036) );
  HS65_LS_NAND2X2 U11595 ( .A(n562), .B(n540), .Z(n6700) );
  HS65_LS_NAND2X2 U11596 ( .A(n36), .B(n14), .Z(n5107) );
  HS65_LS_NAND2X2 U11597 ( .A(n612), .B(n589), .Z(n8152) );
  HS65_LS_NAND2X2 U11598 ( .A(n125), .B(n102), .Z(n8184) );
  HS65_LS_NAND2X2 U11599 ( .A(n837), .B(n826), .Z(n1711) );
  HS65_LS_NAND2X2 U11600 ( .A(n919), .B(n908), .Z(n2463) );
  HS65_LS_NAND2X2 U11601 ( .A(n380), .B(n401), .Z(n7754) );
  HS65_LS_NAND2X2 U11602 ( .A(n217), .B(n204), .Z(n3443) );
  HS65_LS_NAND2X2 U11603 ( .A(n664), .B(n636), .Z(n3687) );
  HS65_LS_NAND2X2 U11604 ( .A(n844), .B(n812), .Z(n1673) );
  HS65_LS_NAND2X2 U11605 ( .A(n926), .B(n894), .Z(n2425) );
  HS65_LS_NAND2X2 U11606 ( .A(n885), .B(n853), .Z(n1297) );
  HS65_LS_NAND2X2 U11607 ( .A(n878), .B(n867), .Z(n1335) );
  HS65_LS_NAND2X2 U11608 ( .A(n803), .B(n771), .Z(n2049) );
  HS65_LS_NAND2X2 U11609 ( .A(n154), .B(n171), .Z(n3587) );
  HS65_LS_NAND2X2 U11610 ( .A(n796), .B(n785), .Z(n2087) );
  HS65_LS_NAND2X2 U11611 ( .A(n640), .B(n656), .Z(n3338) );
  HS65_LS_NAND2X2 U11612 ( .A(n65), .B(n74), .Z(n6849) );
  HS65_LS_NAND2X2 U11613 ( .A(n463), .B(n472), .Z(n5372) );
  HS65_LS_NAND2X2 U11614 ( .A(n286), .B(n295), .Z(n6964) );
  HS65_LS_NAND2X2 U11615 ( .A(n244), .B(n253), .Z(n5257) );
  HS65_LS_NAND2X2 U11616 ( .A(n682), .B(n712), .Z(n5139) );
  HS65_LS_NAND2X2 U11617 ( .A(n500), .B(n530), .Z(n6731) );
  HS65_LS_NAND2X2 U11618 ( .A(n663), .B(n636), .Z(n3172) );
  HS65_LS_NAND2X2 U11619 ( .A(n35), .B(n14), .Z(n4690) );
  HS65_LS_NAND2X2 U11620 ( .A(n561), .B(n540), .Z(n6283) );
  HS65_LS_NAND2X2 U11621 ( .A(n635), .B(n656), .Z(n3713) );
  HS65_LS_NAND2X2 U11622 ( .A(n543), .B(n574), .Z(n6610) );
  HS65_LS_NAND2X2 U11623 ( .A(n17), .B(n48), .Z(n5017) );
  HS65_LS_NAND2X2 U11624 ( .A(n464), .B(n481), .Z(n5408) );
  HS65_LS_NAND2X2 U11625 ( .A(n245), .B(n262), .Z(n5293) );
  HS65_LS_NAND2X2 U11626 ( .A(n680), .B(n700), .Z(n5176) );
  HS65_LS_NAND2X2 U11627 ( .A(n287), .B(n304), .Z(n7000) );
  HS65_LS_NAND2X2 U11628 ( .A(n498), .B(n518), .Z(n6768) );
  HS65_LS_NAND2X2 U11629 ( .A(n66), .B(n83), .Z(n6885) );
  HS65_LS_OAI21X2 U11630 ( .A(n336), .B(n8346), .C(n349), .Z(n8377) );
  HS65_LS_OAI21X2 U11631 ( .A(n547), .B(n548), .C(n566), .Z(n6156) );
  HS65_LS_OAI21X2 U11632 ( .A(n21), .B(n22), .C(n40), .Z(n4563) );
  HS65_LS_NAND2X2 U11633 ( .A(n647), .B(n655), .Z(n3751) );
  HS65_LS_NOR3AX2 U11634 ( .A(n8451), .B(n7985), .C(n8176), .Z(n8437) );
  HS65_LS_NAND2X2 U11635 ( .A(n825), .B(n840), .Z(n1663) );
  HS65_LS_NAND2X2 U11636 ( .A(n907), .B(n922), .Z(n2415) );
  HS65_LS_NAND2X2 U11637 ( .A(n15), .B(n36), .Z(n5054) );
  HS65_LS_NAND2X2 U11638 ( .A(n541), .B(n562), .Z(n6647) );
  HS65_LS_NAND2X2 U11639 ( .A(n639), .B(n660), .Z(n3679) );
  HS65_LS_NOR3AX2 U11640 ( .A(n7866), .B(n8012), .C(n8013), .Z(n7993) );
  HS65_LS_NAND2X2 U11641 ( .A(n784), .B(n799), .Z(n2039) );
  HS65_LS_NAND2X2 U11642 ( .A(n866), .B(n881), .Z(n1287) );
  HS65_LS_NAND2X2 U11643 ( .A(n671), .B(n634), .Z(n3700) );
  HS65_LS_NAND2X2 U11644 ( .A(n192), .B(n228), .Z(n3510) );
  HS65_LS_NOR3AX2 U11645 ( .A(n7949), .B(n8054), .C(n8055), .Z(n8035) );
  HS65_LS_NAND2X2 U11646 ( .A(n440), .B(n413), .Z(n3804) );
  HS65_LS_NAND4ABX3 U11647 ( .A(n2139), .B(n2140), .C(n2141), .D(n2142), .Z(
        n2137) );
  HS65_LS_AOI212X2 U11648 ( .A(n797), .B(n771), .C(n807), .D(n775), .E(n1876), 
        .Z(n2142) );
  HS65_LS_NAND4ABX3 U11649 ( .A(n1387), .B(n1388), .C(n1389), .D(n1390), .Z(
        n1385) );
  HS65_LS_AOI212X2 U11650 ( .A(n879), .B(n853), .C(n889), .D(n857), .E(n1124), 
        .Z(n1390) );
  HS65_LS_OAI21X2 U11651 ( .A(n195), .B(n3085), .C(n227), .Z(n3121) );
  HS65_LS_NAND2X2 U11652 ( .A(n415), .B(n436), .Z(n3796) );
  HS65_LS_NAND2X2 U11653 ( .A(n199), .B(n214), .Z(n3435) );
  HS65_LS_NAND2X2 U11654 ( .A(n423), .B(n431), .Z(n3868) );
  HS65_LS_NAND2X2 U11655 ( .A(n336), .B(n353), .Z(n8617) );
  HS65_LS_OAI21X2 U11656 ( .A(n373), .B(n8093), .C(n390), .Z(n8092) );
  HS65_LS_NAND2X2 U11657 ( .A(n352), .B(n326), .Z(n8050) );
  HS65_LS_NAND2X2 U11658 ( .A(n643), .B(n663), .Z(n3688) );
  HS65_LS_NAND2X2 U11659 ( .A(n331), .B(n344), .Z(n7771) );
  HS65_LS_NAND2X2 U11660 ( .A(n191), .B(n213), .Z(n3439) );
  HS65_LS_NAND2X2 U11661 ( .A(n16), .B(n48), .Z(n5044) );
  HS65_LS_NAND2X2 U11662 ( .A(n542), .B(n574), .Z(n6637) );
  HS65_LS_NAND2X2 U11663 ( .A(n542), .B(n562), .Z(n6678) );
  HS65_LS_NAND2X2 U11664 ( .A(n16), .B(n36), .Z(n5085) );
  HS65_LS_NAND2X2 U11665 ( .A(n217), .B(n193), .Z(n3110) );
  HS65_LS_OAI21X2 U11666 ( .A(n199), .B(n3085), .C(n223), .Z(n3904) );
  HS65_LS_NOR3X1 U11667 ( .A(n7910), .B(n7658), .C(n7728), .Z(n7876) );
  HS65_LS_NAND2X2 U11668 ( .A(n920), .B(n904), .Z(n2444) );
  HS65_LS_NAND2X2 U11669 ( .A(n838), .B(n822), .Z(n1692) );
  HS65_LS_OAI21X2 U11670 ( .A(n329), .B(n8346), .C(n354), .Z(n8882) );
  HS65_LS_NAND2X2 U11671 ( .A(n378), .B(n401), .Z(n8233) );
  HS65_LS_NAND2X2 U11672 ( .A(n646), .B(n663), .Z(n3746) );
  HS65_LS_NAND2X2 U11673 ( .A(n879), .B(n863), .Z(n1316) );
  HS65_LS_NAND2X2 U11674 ( .A(n797), .B(n781), .Z(n2068) );
  HS65_LS_NAND2X2 U11675 ( .A(n56), .B(n80), .Z(n6949) );
  HS65_LS_NAND2X2 U11676 ( .A(n454), .B(n478), .Z(n5472) );
  HS65_LS_NAND2X2 U11677 ( .A(n277), .B(n301), .Z(n7064) );
  HS65_LS_NAND2X2 U11678 ( .A(n235), .B(n259), .Z(n5357) );
  HS65_LS_NAND2X2 U11679 ( .A(n688), .B(n697), .Z(n5242) );
  HS65_LS_NAND2X2 U11680 ( .A(n506), .B(n515), .Z(n6834) );
  HS65_LS_NAND2X2 U11681 ( .A(n462), .B(n472), .Z(n5398) );
  HS65_LS_NAND2X2 U11682 ( .A(n243), .B(n253), .Z(n5283) );
  HS65_LS_NAND2X2 U11683 ( .A(n285), .B(n295), .Z(n6990) );
  HS65_LS_NAND2X2 U11684 ( .A(n681), .B(n712), .Z(n5166) );
  HS65_LS_NAND2X2 U11685 ( .A(n64), .B(n74), .Z(n6875) );
  HS65_LS_NAND2X2 U11686 ( .A(n499), .B(n530), .Z(n6758) );
  HS65_LS_NAND2X2 U11687 ( .A(n583), .B(n615), .Z(n7807) );
  HS65_LS_NAND2X2 U11688 ( .A(n96), .B(n128), .Z(n7907) );
  HS65_LS_NAND2X2 U11689 ( .A(n925), .B(n894), .Z(n2380) );
  HS65_LS_NAND2X2 U11690 ( .A(n843), .B(n812), .Z(n1628) );
  HS65_LS_NAND2X2 U11691 ( .A(n649), .B(n659), .Z(n3684) );
  HS65_LS_NAND2X2 U11692 ( .A(n76), .B(n60), .Z(n6915) );
  HS65_LS_NAND2X2 U11693 ( .A(n255), .B(n239), .Z(n5323) );
  HS65_LS_NAND2X2 U11694 ( .A(n474), .B(n458), .Z(n5438) );
  HS65_LS_NAND2X2 U11695 ( .A(n297), .B(n281), .Z(n7030) );
  HS65_LS_NAND2X2 U11696 ( .A(n710), .B(n683), .Z(n5207) );
  HS65_LS_NAND2X2 U11697 ( .A(n528), .B(n501), .Z(n6799) );
  HS65_LS_NAND2X2 U11698 ( .A(n909), .B(n928), .Z(n2363) );
  HS65_LS_NAND2X2 U11699 ( .A(n827), .B(n846), .Z(n1611) );
  HS65_LS_NAND2X2 U11700 ( .A(n884), .B(n853), .Z(n1252) );
  HS65_LS_NAND2X2 U11701 ( .A(n550), .B(n559), .Z(n6699) );
  HS65_LS_NAND2X2 U11702 ( .A(n24), .B(n33), .Z(n5106) );
  HS65_LS_NAND2X2 U11703 ( .A(n419), .B(n435), .Z(n3849) );
  HS65_LS_NAND2X2 U11704 ( .A(n379), .B(n397), .Z(n8090) );
  HS65_LS_NAND2X2 U11705 ( .A(n868), .B(n887), .Z(n1235) );
  HS65_LS_NAND2X2 U11706 ( .A(n786), .B(n805), .Z(n1987) );
  HS65_LS_NAND2X2 U11707 ( .A(n802), .B(n771), .Z(n2004) );
  HS65_LS_NOR3AX2 U11708 ( .A(n6492), .B(n6332), .C(n6190), .Z(n6475) );
  HS65_LS_NOR3AX2 U11709 ( .A(n4682), .B(n4554), .C(n4483), .Z(n4664) );
  HS65_LS_NOR3AX2 U11710 ( .A(n6275), .B(n6147), .C(n6076), .Z(n6257) );
  HS65_LS_NOR3AX2 U11711 ( .A(n4899), .B(n4739), .C(n4597), .Z(n4882) );
  HS65_LS_NAND2X2 U11712 ( .A(n903), .B(n926), .Z(n2431) );
  HS65_LS_NAND2X2 U11713 ( .A(n821), .B(n844), .Z(n1679) );
  HS65_LS_NAND2X2 U11714 ( .A(n168), .B(n159), .Z(n3657) );
  HS65_LS_NAND2X2 U11715 ( .A(n586), .B(n618), .Z(n8710) );
  HS65_LS_NAND2X2 U11716 ( .A(n99), .B(n131), .Z(n8798) );
  HS65_LS_NAND2X2 U11717 ( .A(n543), .B(n568), .Z(n6648) );
  HS65_LS_NAND2X2 U11718 ( .A(n17), .B(n42), .Z(n5055) );
  HS65_LS_NAND2X2 U11719 ( .A(n639), .B(n670), .Z(n3358) );
  HS65_LS_NAND2X2 U11720 ( .A(n862), .B(n885), .Z(n1303) );
  HS65_LS_NAND2X2 U11721 ( .A(n780), .B(n803), .Z(n2055) );
  HS65_LS_NAND2X2 U11722 ( .A(n571), .B(n537), .Z(n6083) );
  HS65_LS_NAND2X2 U11723 ( .A(n45), .B(n11), .Z(n4490) );
  HS65_LS_NAND2X2 U11724 ( .A(n327), .B(n350), .Z(n8354) );
  HS65_LS_NAND2X2 U11725 ( .A(n709), .B(n676), .Z(n4546) );
  HS65_LS_NAND2X2 U11726 ( .A(n475), .B(n468), .Z(n4615) );
  HS65_LS_NAND2X2 U11727 ( .A(n298), .B(n291), .Z(n6208) );
  HS65_LS_NAND2X2 U11728 ( .A(n77), .B(n70), .Z(n6196) );
  HS65_LS_NAND2X2 U11729 ( .A(n527), .B(n494), .Z(n6139) );
  HS65_LS_NAND2X2 U11730 ( .A(n256), .B(n249), .Z(n4603) );
  HS65_LS_NAND2X2 U11731 ( .A(n667), .B(n635), .Z(n3760) );
  HS65_LS_NAND2X2 U11732 ( .A(n917), .B(n904), .Z(n2412) );
  HS65_LS_NAND2X2 U11733 ( .A(n835), .B(n822), .Z(n1660) );
  HS65_LS_OAI21X2 U11734 ( .A(n639), .B(n3314), .C(n669), .Z(n3965) );
  HS65_LS_NAND2X2 U11735 ( .A(n439), .B(n412), .Z(n3836) );
  HS65_LS_NAND4ABX3 U11736 ( .A(n3612), .B(n3613), .C(n3614), .D(n3615), .Z(
        n3028) );
  HS65_LS_NOR3X1 U11737 ( .A(n3620), .B(n3621), .C(n3622), .Z(n3614) );
  HS65_LS_NOR4ABX2 U11738 ( .A(n3616), .B(n3617), .C(n3618), .D(n3619), .Z(
        n3615) );
  HS65_LS_NAND4ABX3 U11739 ( .A(n3626), .B(n3627), .C(n3628), .D(n3629), .Z(
        n3612) );
  HS65_LS_NAND2X2 U11740 ( .A(n876), .B(n863), .Z(n1284) );
  HS65_LS_NAND2X2 U11741 ( .A(n794), .B(n781), .Z(n2036) );
  HS65_LS_NAND2X2 U11742 ( .A(n345), .B(n336), .Z(n8353) );
  HS65_LS_OAI21X2 U11743 ( .A(n378), .B(n8093), .C(n391), .Z(n8508) );
  HS65_LS_NAND2X2 U11744 ( .A(n381), .B(n390), .Z(n8240) );
  HS65_LS_NAND2X2 U11745 ( .A(n437), .B(n421), .Z(n3383) );
  HS65_LS_NAND2X2 U11746 ( .A(n439), .B(n421), .Z(n3400) );
  HS65_LS_NAND4ABX3 U11747 ( .A(n8558), .B(n8559), .C(n8560), .D(n8561), .Z(
        n8053) );
  HS65_LS_NOR3AX2 U11748 ( .A(n8566), .B(n8567), .C(n8568), .Z(n8560) );
  HS65_LS_NAND4ABX3 U11749 ( .A(n8572), .B(n8573), .C(n7771), .D(n8574), .Z(
        n8558) );
  HS65_LS_NOR4ABX2 U11750 ( .A(n8562), .B(n8563), .C(n8564), .D(n8565), .Z(
        n8561) );
  HS65_LS_NAND2X2 U11751 ( .A(n199), .B(n221), .Z(n3132) );
  HS65_LS_NAND2X2 U11752 ( .A(n415), .B(n446), .Z(n3420) );
  HS65_LS_NAND4ABX3 U11753 ( .A(n3714), .B(n3715), .C(n3716), .D(n3717), .Z(
        n3139) );
  HS65_LS_NAND4ABX3 U11754 ( .A(n3729), .B(n3730), .C(n3731), .D(n3732), .Z(
        n3714) );
  HS65_LS_NOR4ABX2 U11755 ( .A(n3718), .B(n3719), .C(n3720), .D(n3721), .Z(
        n3717) );
  HS65_LS_NOR3AX2 U11756 ( .A(n3722), .B(n3723), .C(n3724), .Z(n3716) );
  HS65_LS_NAND2X2 U11757 ( .A(n425), .B(n435), .Z(n3801) );
  HS65_LS_NAND4ABX3 U11758 ( .A(n3472), .B(n3473), .C(n3474), .D(n3475), .Z(
        n2936) );
  HS65_LS_NOR3X1 U11759 ( .A(n3480), .B(n3481), .C(n3482), .Z(n3474) );
  HS65_LS_NAND4ABX3 U11760 ( .A(n3487), .B(n3488), .C(n3489), .D(n3490), .Z(
        n3472) );
  HS65_LS_NOR4ABX2 U11761 ( .A(n3476), .B(n3477), .C(n3478), .D(n3479), .Z(
        n3475) );
  HS65_LS_NAND2X2 U11762 ( .A(n148), .B(n176), .Z(n3035) );
  HS65_LS_NAND4ABX3 U11763 ( .A(n8254), .B(n8255), .C(n8256), .D(n8257), .Z(
        n8011) );
  HS65_LS_NOR3AX2 U11764 ( .A(n8262), .B(n8263), .C(n8264), .Z(n8256) );
  HS65_LS_NAND4ABX3 U11765 ( .A(n8268), .B(n8269), .C(n8270), .D(n7754), .Z(
        n8254) );
  HS65_LS_NOR4ABX2 U11766 ( .A(n8258), .B(n8259), .C(n8260), .D(n8261), .Z(
        n8257) );
  HS65_LS_NAND2X2 U11767 ( .A(n127), .B(n110), .Z(n7904) );
  HS65_LS_NAND2X2 U11768 ( .A(n614), .B(n597), .Z(n7804) );
  HS65_LS_NAND2X2 U11769 ( .A(n172), .B(n159), .Z(n3566) );
  HS65_LS_NAND2X2 U11770 ( .A(n583), .B(n609), .Z(n8703) );
  HS65_LS_NAND2X2 U11771 ( .A(n96), .B(n122), .Z(n8791) );
  HS65_LS_NAND2X2 U11772 ( .A(n661), .B(n645), .Z(n3321) );
  HS65_LS_NOR3AX2 U11773 ( .A(n3366), .B(n3378), .C(n3180), .Z(n3819) );
  HS65_LS_NAND2X2 U11774 ( .A(n640), .B(n665), .Z(n3151) );
  HS65_LS_NAND2X2 U11775 ( .A(n201), .B(n216), .Z(n2949) );
  HS65_LS_NAND2X2 U11776 ( .A(n416), .B(n441), .Z(n3192) );
  HS65_LS_NAND2X2 U11777 ( .A(n404), .B(n373), .Z(n8111) );
  HS65_LS_NAND2X2 U11778 ( .A(n58), .B(n88), .Z(n6934) );
  HS65_LS_NAND2X2 U11779 ( .A(n237), .B(n267), .Z(n5342) );
  HS65_LS_NAND2X2 U11780 ( .A(n456), .B(n486), .Z(n5457) );
  HS65_LS_NAND2X2 U11781 ( .A(n279), .B(n309), .Z(n7049) );
  HS65_LS_NAND2X2 U11782 ( .A(n508), .B(n523), .Z(n6818) );
  HS65_LS_NAND2X2 U11783 ( .A(n690), .B(n705), .Z(n5226) );
  HS65_LS_NAND2X2 U11784 ( .A(n552), .B(n567), .Z(n6713) );
  HS65_LS_NAND2X2 U11785 ( .A(n26), .B(n41), .Z(n5120) );
  HS65_LS_NAND2X2 U11786 ( .A(n218), .B(n202), .Z(n3477) );
  HS65_LS_NAND2X2 U11787 ( .A(n366), .B(n394), .Z(n8120) );
  HS65_LS_NAND2X2 U11788 ( .A(n354), .B(n336), .Z(n8584) );
  HS65_LS_NAND2X2 U11789 ( .A(n372), .B(n399), .Z(n8279) );
  HS65_LS_NAND2X2 U11790 ( .A(n445), .B(n421), .Z(n3864) );
  HS65_LS_NAND2X2 U11791 ( .A(n548), .B(n567), .Z(n6305) );
  HS65_LS_NAND2X2 U11792 ( .A(n22), .B(n41), .Z(n4712) );
  HS65_LS_NAND2X2 U11793 ( .A(n170), .B(n150), .Z(n3561) );
  HS65_LS_NAND2X2 U11794 ( .A(n593), .B(n615), .Z(n8721) );
  HS65_LS_NAND2X2 U11795 ( .A(n106), .B(n128), .Z(n8809) );
  HS65_LS_NAND2X2 U11796 ( .A(n586), .B(n615), .Z(n8417) );
  HS65_LS_NAND2X2 U11797 ( .A(n99), .B(n128), .Z(n8477) );
  HS65_LS_NAND2X2 U11798 ( .A(n110), .B(n138), .Z(n7920) );
  HS65_LS_NAND2X2 U11799 ( .A(n597), .B(n625), .Z(n7821) );
  HS65_LS_NAND2X2 U11800 ( .A(n643), .B(n659), .Z(n3731) );
  HS65_LS_NAND4ABX3 U11801 ( .A(n8691), .B(n8692), .C(n8693), .D(n8694), .Z(
        n8142) );
  HS65_LS_NAND4ABX3 U11802 ( .A(n7820), .B(n8702), .C(n8703), .D(n7680), .Z(
        n8691) );
  HS65_LS_NOR4ABX2 U11803 ( .A(n8695), .B(n8696), .C(n7707), .D(n7799), .Z(
        n8694) );
  HS65_LS_NOR3AX2 U11804 ( .A(n8697), .B(n7840), .C(n8698), .Z(n8693) );
  HS65_LS_NAND4ABX3 U11805 ( .A(n8779), .B(n8780), .C(n8781), .D(n8782), .Z(
        n8174) );
  HS65_LS_NAND4ABX3 U11806 ( .A(n7919), .B(n8790), .C(n8791), .D(n7718), .Z(
        n8779) );
  HS65_LS_NOR4ABX2 U11807 ( .A(n8783), .B(n8784), .C(n7745), .D(n7899), .Z(
        n8782) );
  HS65_LS_NOR3AX2 U11808 ( .A(n8785), .B(n7939), .C(n8786), .Z(n8781) );
  HS65_LS_NAND2X2 U11809 ( .A(n154), .B(n175), .Z(n3296) );
  HS65_LS_NAND2X2 U11810 ( .A(n327), .B(n346), .Z(n8570) );
  HS65_LS_NAND2X2 U11811 ( .A(n64), .B(n83), .Z(n6914) );
  HS65_LS_NAND2X2 U11812 ( .A(n243), .B(n262), .Z(n5322) );
  HS65_LS_NAND2X2 U11813 ( .A(n462), .B(n481), .Z(n5437) );
  HS65_LS_NAND2X2 U11814 ( .A(n285), .B(n304), .Z(n7029) );
  HS65_LS_NAND2X2 U11815 ( .A(n681), .B(n700), .Z(n5206) );
  HS65_LS_NAND2X2 U11816 ( .A(n499), .B(n518), .Z(n6798) );
  HS65_LS_NAND2X2 U11817 ( .A(n167), .B(n150), .Z(n3583) );
  HS65_LS_NAND2X2 U11818 ( .A(n391), .B(n373), .Z(n8280) );
  HS65_LS_NAND2X2 U11819 ( .A(n901), .B(n926), .Z(n2472) );
  HS65_LS_NAND2X2 U11820 ( .A(n819), .B(n844), .Z(n1720) );
  HS65_LS_NAND2X2 U11821 ( .A(n193), .B(n213), .Z(n3489) );
  HS65_LS_NAND2X2 U11822 ( .A(n56), .B(n88), .Z(n6486) );
  HS65_LS_NAND2X2 U11823 ( .A(n277), .B(n309), .Z(n6600) );
  HS65_LS_NAND2X2 U11824 ( .A(n235), .B(n267), .Z(n4893) );
  HS65_LS_NAND2X2 U11825 ( .A(n454), .B(n486), .Z(n5007) );
  HS65_LS_NAND2X2 U11826 ( .A(n688), .B(n705), .Z(n4879) );
  HS65_LS_NAND2X2 U11827 ( .A(n506), .B(n523), .Z(n6472) );
  HS65_LS_NAND2X2 U11828 ( .A(n24), .B(n41), .Z(n4675) );
  HS65_LS_NAND2X2 U11829 ( .A(n550), .B(n567), .Z(n6268) );
  HS65_LS_OAI21X2 U11830 ( .A(n421), .B(n3376), .C(n430), .Z(n3410) );
  HS65_LS_NAND2X2 U11831 ( .A(n860), .B(n885), .Z(n1344) );
  HS65_LS_NAND2X2 U11832 ( .A(n778), .B(n803), .Z(n2096) );
  HS65_LS_NAND2X2 U11833 ( .A(n212), .B(n195), .Z(n3092) );
  HS65_LS_NAND2X2 U11834 ( .A(n218), .B(n195), .Z(n3111) );
  HS65_LS_NAND2X2 U11835 ( .A(n925), .B(n900), .Z(n2304) );
  HS65_LS_NAND2X2 U11836 ( .A(n843), .B(n818), .Z(n1552) );
  HS65_LS_NAND2X2 U11837 ( .A(n16), .B(n32), .Z(n5058) );
  HS65_LS_NAND2X2 U11838 ( .A(n542), .B(n558), .Z(n6651) );
  HS65_LS_NAND2X2 U11839 ( .A(n650), .B(n670), .Z(n3331) );
  HS65_LS_NAND2X2 U11840 ( .A(n374), .B(n399), .Z(n8259) );
  HS65_LS_NAND2X2 U11841 ( .A(n598), .B(n625), .Z(n8434) );
  HS65_LS_NAND2X2 U11842 ( .A(n111), .B(n138), .Z(n8445) );
  HS65_LS_NAND2X2 U11843 ( .A(n443), .B(n412), .Z(n3877) );
  HS65_LS_NAND2X2 U11844 ( .A(n608), .B(n599), .Z(n8731) );
  HS65_LS_NAND2X2 U11845 ( .A(n121), .B(n112), .Z(n8819) );
  HS65_LS_NAND2X2 U11846 ( .A(n884), .B(n859), .Z(n1176) );
  HS65_LS_OAI21X2 U11847 ( .A(n177), .B(n3050), .C(n158), .Z(n3049) );
  HS65_LS_NAND2X2 U11848 ( .A(n596), .B(n615), .Z(n8397) );
  HS65_LS_NAND2X2 U11849 ( .A(n109), .B(n128), .Z(n8457) );
  HS65_LS_NAND2X2 U11850 ( .A(n62), .B(n88), .Z(n6521) );
  HS65_LS_NAND2X2 U11851 ( .A(n460), .B(n486), .Z(n4982) );
  HS65_LS_NAND2X2 U11852 ( .A(n283), .B(n309), .Z(n6575) );
  HS65_LS_NAND2X2 U11853 ( .A(n241), .B(n267), .Z(n4928) );
  HS65_LS_NAND2X2 U11854 ( .A(n686), .B(n705), .Z(n4852) );
  HS65_LS_NAND2X2 U11855 ( .A(n504), .B(n523), .Z(n6445) );
  HS65_LS_NAND2X2 U11856 ( .A(n802), .B(n777), .Z(n1928) );
  HS65_LS_NAND2X2 U11857 ( .A(n22), .B(n48), .Z(n5040) );
  HS65_LS_NAND2X2 U11858 ( .A(n548), .B(n574), .Z(n6633) );
  HS65_LS_NAND2X2 U11859 ( .A(n323), .B(n352), .Z(n8376) );
  HS65_LS_NAND2X2 U11860 ( .A(n903), .B(n928), .Z(n2379) );
  HS65_LS_NAND2X2 U11861 ( .A(n821), .B(n846), .Z(n1627) );
  HS65_LS_OAI21X2 U11862 ( .A(n415), .B(n3376), .C(n445), .Z(n3986) );
  HS65_LS_NAND2X2 U11863 ( .A(n930), .B(n910), .Z(n2373) );
  HS65_LS_NAND2X2 U11864 ( .A(n848), .B(n828), .Z(n1621) );
  HS65_LS_NAND2X2 U11865 ( .A(n807), .B(n787), .Z(n1997) );
  HS65_LS_NAND2X2 U11866 ( .A(n889), .B(n869), .Z(n1245) );
  HS65_LS_NAND2X2 U11867 ( .A(n862), .B(n887), .Z(n1251) );
  HS65_LS_NAND2X2 U11868 ( .A(n780), .B(n805), .Z(n2003) );
  HS65_LS_NAND2X2 U11869 ( .A(n462), .B(n477), .Z(n5412) );
  HS65_LS_NAND2X2 U11870 ( .A(n243), .B(n258), .Z(n5297) );
  HS65_LS_NAND2X2 U11871 ( .A(n285), .B(n300), .Z(n7004) );
  HS65_LS_NAND2X2 U11872 ( .A(n681), .B(n696), .Z(n5180) );
  HS65_LS_NAND2X2 U11873 ( .A(n499), .B(n514), .Z(n6772) );
  HS65_LS_NAND2X2 U11874 ( .A(n64), .B(n79), .Z(n6889) );
  HS65_LS_NAND2X2 U11875 ( .A(n426), .B(n446), .Z(n3393) );
  HS65_LS_NAND2X2 U11876 ( .A(n190), .B(n221), .Z(n3104) );
  HS65_LS_NAND2X2 U11877 ( .A(n585), .B(n618), .Z(n7800) );
  HS65_LS_NAND2X2 U11878 ( .A(n98), .B(n131), .Z(n7900) );
  HS65_LS_NAND2X2 U11879 ( .A(n199), .B(n222), .Z(n3440) );
  HS65_LS_NAND2X2 U11880 ( .A(n223), .B(n195), .Z(n3506) );
  HS65_LS_NAND2X2 U11881 ( .A(n219), .B(n202), .Z(n3519) );
  HS65_LS_NAND2X2 U11882 ( .A(n352), .B(n336), .Z(n8369) );
  HS65_LS_NAND2X2 U11883 ( .A(n180), .B(n157), .Z(n3606) );
  HS65_LS_NAND2X2 U11884 ( .A(n156), .B(n175), .Z(n3582) );
  HS65_LS_OAI21X2 U11885 ( .A(n193), .B(n189), .C(n212), .Z(n4235) );
  HS65_LS_NAND2X2 U11886 ( .A(n670), .B(n644), .Z(n3709) );
  HS65_LS_NOR3AX2 U11887 ( .A(n3286), .B(n3287), .C(n3288), .Z(n3274) );
  HS65_LS_OAI21X2 U11888 ( .A(n150), .B(n3247), .C(n181), .Z(n3286) );
  HS65_LS_NAND2X2 U11889 ( .A(n176), .B(n159), .Z(n3656) );
  HS65_LS_NAND2X2 U11890 ( .A(n663), .B(n645), .Z(n3337) );
  HS65_LS_NAND2X2 U11891 ( .A(n394), .B(n371), .Z(n8248) );
  HS65_LS_NAND2X2 U11892 ( .A(n177), .B(n150), .Z(n3258) );
  HS65_LS_NAND2X2 U11893 ( .A(n399), .B(n373), .Z(n8127) );
  HS65_LS_NAND2X2 U11894 ( .A(n649), .B(n658), .Z(n3737) );
  HS65_LS_NAND4ABX3 U11895 ( .A(n6075), .B(n6076), .C(n6077), .D(n6078), .Z(
        n6074) );
  HS65_LS_AOI212X2 U11896 ( .A(n541), .B(n559), .C(n537), .D(n574), .E(n6079), 
        .Z(n6078) );
  HS65_LS_NAND4ABX3 U11897 ( .A(n4482), .B(n4483), .C(n4484), .D(n4485), .Z(
        n4481) );
  HS65_LS_AOI212X2 U11898 ( .A(n15), .B(n33), .C(n11), .D(n48), .E(n4486), .Z(
        n4485) );
  HS65_LS_NAND4ABX3 U11899 ( .A(n4608), .B(n4609), .C(n4610), .D(n4611), .Z(
        n4607) );
  HS65_LS_AOI212X2 U11900 ( .A(n464), .B(n478), .C(n468), .D(n472), .E(n4612), 
        .Z(n4611) );
  HS65_LS_NAND4ABX3 U11901 ( .A(n6201), .B(n6202), .C(n6203), .D(n6204), .Z(
        n6200) );
  HS65_LS_AOI212X2 U11902 ( .A(n287), .B(n301), .C(n291), .D(n295), .E(n6205), 
        .Z(n6204) );
  HS65_LS_NAND2X2 U11903 ( .A(n221), .B(n197), .Z(n3466) );
  HS65_LS_NAND2X2 U11904 ( .A(n917), .B(n905), .Z(n2449) );
  HS65_LS_NAND2X2 U11905 ( .A(n835), .B(n823), .Z(n1697) );
  HS65_LS_NAND2X2 U11906 ( .A(n542), .B(n567), .Z(n6677) );
  HS65_LS_NAND2X2 U11907 ( .A(n16), .B(n41), .Z(n5084) );
  HS65_LS_OAI21X2 U11908 ( .A(n148), .B(n143), .C(n166), .Z(n4173) );
  HS65_LS_NAND2X2 U11909 ( .A(n42), .B(n22), .Z(n5079) );
  HS65_LS_NAND2X2 U11910 ( .A(n568), .B(n548), .Z(n6672) );
  HS65_LS_NAND2X2 U11911 ( .A(n356), .B(n337), .Z(n8552) );
  HS65_LS_NAND2X2 U11912 ( .A(n876), .B(n864), .Z(n1321) );
  HS65_LS_NAND2X2 U11913 ( .A(n794), .B(n782), .Z(n2073) );
  HS65_LS_NAND2X2 U11914 ( .A(n425), .B(n434), .Z(n3854) );
  HS65_LS_NAND2X2 U11915 ( .A(n321), .B(n348), .Z(n7966) );
  HS65_LS_NAND2X2 U11916 ( .A(n176), .B(n150), .Z(n3648) );
  HS65_LS_NAND4ABX3 U11917 ( .A(n7971), .B(n7972), .C(n7973), .D(n7974), .Z(
        n7970) );
  HS65_LS_AOI212X2 U11918 ( .A(n622), .B(n584), .C(n592), .D(n609), .E(n7975), 
        .Z(n7974) );
  HS65_LS_NAND4ABX3 U11919 ( .A(n7984), .B(n7985), .C(n7986), .D(n7987), .Z(
        n7983) );
  HS65_LS_AOI212X2 U11920 ( .A(n135), .B(n97), .C(n105), .D(n122), .E(n7988), 
        .Z(n7987) );
  HS65_LS_OAI21X2 U11921 ( .A(n594), .B(n8400), .C(n618), .Z(n9062) );
  HS65_LS_OAI21X2 U11922 ( .A(n107), .B(n8460), .C(n131), .Z(n9120) );
  HS65_LS_OAI21X2 U11923 ( .A(n354), .B(n353), .C(n321), .Z(n8905) );
  HS65_LS_NAND2X2 U11924 ( .A(n650), .B(n658), .Z(n2991) );
  HS65_LS_OAI21X2 U11925 ( .A(n818), .B(n822), .C(n836), .Z(n1842) );
  HS65_LS_OAI21X2 U11926 ( .A(n900), .B(n904), .C(n918), .Z(n2594) );
  HS65_LS_NAND2X2 U11927 ( .A(n366), .B(n388), .Z(n7864) );
  HS65_LS_NAND2X2 U11928 ( .A(n930), .B(n905), .Z(n2288) );
  HS65_LS_NAND2X2 U11929 ( .A(n848), .B(n823), .Z(n1536) );
  HS65_LS_OAI21X2 U11930 ( .A(n391), .B(n396), .C(n366), .Z(n8965) );
  HS65_LS_NAND2X2 U11931 ( .A(n377), .B(n386), .Z(n8258) );
  HS65_LS_OAI21X2 U11932 ( .A(n777), .B(n781), .C(n795), .Z(n2218) );
  HS65_LS_OAI21X2 U11933 ( .A(n859), .B(n863), .C(n877), .Z(n1466) );
  HS65_LS_NAND2X2 U11934 ( .A(n191), .B(n225), .Z(n3495) );
  HS65_LS_NAND2X2 U11935 ( .A(n889), .B(n864), .Z(n1160) );
  HS65_LS_NAND2X2 U11936 ( .A(n807), .B(n782), .Z(n1912) );
  HS65_LS_OAI21X2 U11937 ( .A(n160), .B(n143), .C(n171), .Z(n3279) );
  HS65_LS_OAI21X2 U11938 ( .A(n901), .B(n899), .C(n928), .Z(n2337) );
  HS65_LS_OAI21X2 U11939 ( .A(n819), .B(n817), .C(n846), .Z(n1585) );
  HS65_LS_NAND2X2 U11940 ( .A(n426), .B(n434), .Z(n3009) );
  HS65_LS_NAND2X2 U11941 ( .A(n404), .B(n371), .Z(n8302) );
  HS65_LS_OAI21X2 U11942 ( .A(n65), .B(n63), .C(n77), .Z(n7475) );
  HS65_LS_OAI21X2 U11943 ( .A(n463), .B(n461), .C(n475), .Z(n5942) );
  HS65_LS_OAI21X2 U11944 ( .A(n286), .B(n284), .C(n298), .Z(n7534) );
  HS65_LS_OAI21X2 U11945 ( .A(n244), .B(n242), .C(n256), .Z(n5883) );
  HS65_LS_OAI21X2 U11946 ( .A(n682), .B(n679), .C(n709), .Z(n5776) );
  HS65_LS_OAI21X2 U11947 ( .A(n500), .B(n497), .C(n527), .Z(n7368) );
  HS65_LS_OAI21X2 U11948 ( .A(n35), .B(n43), .C(n20), .Z(n5759) );
  HS65_LS_OAI21X2 U11949 ( .A(n561), .B(n569), .C(n546), .Z(n7351) );
  HS65_LS_OAI21X2 U11950 ( .A(n667), .B(n665), .C(n644), .Z(n4029) );
  HS65_LS_OAI21X2 U11951 ( .A(n860), .B(n858), .C(n887), .Z(n1209) );
  HS65_LS_OAI21X2 U11952 ( .A(n778), .B(n776), .C(n805), .Z(n1961) );
  HS65_LS_NAND2X2 U11953 ( .A(n589), .B(n611), .Z(n8418) );
  HS65_LS_NAND2X2 U11954 ( .A(n102), .B(n124), .Z(n8478) );
  HS65_LS_OAI21X2 U11955 ( .A(n89), .B(n85), .C(n64), .Z(n7212) );
  HS65_LS_OAI21X2 U11956 ( .A(n487), .B(n483), .C(n462), .Z(n5647) );
  HS65_LS_OAI21X2 U11957 ( .A(n310), .B(n306), .C(n285), .Z(n7239) );
  HS65_LS_OAI21X2 U11958 ( .A(n268), .B(n264), .C(n243), .Z(n5620) );
  HS65_LS_OAI21X2 U11959 ( .A(n704), .B(n701), .C(n681), .Z(n5593) );
  HS65_LS_OAI21X2 U11960 ( .A(n522), .B(n519), .C(n499), .Z(n7185) );
  HS65_LS_OAI21X2 U11961 ( .A(n773), .B(n774), .C(n792), .Z(n2154) );
  HS65_LS_OAI21X2 U11962 ( .A(n855), .B(n856), .C(n874), .Z(n1402) );
  HS65_LS_OAI21X2 U11963 ( .A(n814), .B(n815), .C(n833), .Z(n1778) );
  HS65_LS_OAI21X2 U11964 ( .A(n896), .B(n897), .C(n915), .Z(n2530) );
  HS65_LS_OAI21X2 U11965 ( .A(n169), .B(n177), .C(n158), .Z(n4166) );
  HS65_LS_OAI21X2 U11966 ( .A(n543), .B(n540), .C(n571), .Z(n7306) );
  HS65_LS_OAI21X2 U11967 ( .A(n17), .B(n14), .C(n45), .Z(n5714) );
  HS65_LS_NAND2X2 U11968 ( .A(n331), .B(n348), .Z(n8579) );
  HS65_LS_NAND2X2 U11969 ( .A(n35), .B(n16), .Z(n5103) );
  HS65_LS_NAND2X2 U11970 ( .A(n561), .B(n542), .Z(n6696) );
  HS65_LS_OAI21X2 U11971 ( .A(n215), .B(n222), .C(n203), .Z(n4200) );
  HS65_LS_OAI21X2 U11972 ( .A(n219), .B(n216), .C(n197), .Z(n3944) );
  HS65_LS_OAI21X2 U11973 ( .A(n443), .B(n441), .C(n420), .Z(n4053) );
  HS65_LS_NOR3AX2 U11974 ( .A(n3199), .B(n3200), .C(n3201), .Z(n3183) );
  HS65_LS_OAI21X2 U11975 ( .A(n174), .B(n168), .C(n150), .Z(n3291) );
  HS65_LS_OAI21X2 U11976 ( .A(n350), .B(n358), .C(n323), .Z(n8873) );
  HS65_LS_NAND2X2 U11977 ( .A(n655), .B(n644), .Z(n3718) );
  HS65_LS_OAI21X2 U11978 ( .A(n484), .B(n4523), .C(n458), .Z(n4521) );
  HS65_LS_OAI21X2 U11979 ( .A(n265), .B(n4477), .C(n239), .Z(n4475) );
  HS65_LS_OAI21X2 U11980 ( .A(n307), .B(n6116), .C(n281), .Z(n6114) );
  HS65_LS_OAI21X2 U11981 ( .A(n699), .B(n5505), .C(n683), .Z(n5827) );
  HS65_LS_OAI21X2 U11982 ( .A(n35), .B(n5489), .C(n18), .Z(n5765) );
  HS65_LS_OAI21X2 U11983 ( .A(n517), .B(n7097), .C(n501), .Z(n7419) );
  HS65_LS_OAI21X2 U11984 ( .A(n86), .B(n6070), .C(n60), .Z(n6068) );
  HS65_LS_OAI21X2 U11985 ( .A(n561), .B(n7081), .C(n544), .Z(n7357) );
  HS65_LS_OAI21X2 U11986 ( .A(n616), .B(n622), .C(n586), .Z(n8431) );
  HS65_LS_OAI21X2 U11987 ( .A(n129), .B(n135), .C(n99), .Z(n8442) );
  HS65_LS_OAI21X2 U11988 ( .A(n174), .B(n170), .C(n152), .Z(n4005) );
  HS65_LS_OAI21X2 U11989 ( .A(n612), .B(n620), .C(n600), .Z(n9031) );
  HS65_LS_OAI21X2 U11990 ( .A(n125), .B(n133), .C(n113), .Z(n9089) );
  HS65_LS_OAI21X2 U11991 ( .A(n895), .B(n910), .C(n923), .Z(n2285) );
  HS65_LS_OAI21X2 U11992 ( .A(n813), .B(n828), .C(n841), .Z(n1533) );
  HS65_LS_OAI21X2 U11993 ( .A(n613), .B(n623), .C(n599), .Z(n8435) );
  HS65_LS_NAND2X2 U11994 ( .A(n484), .B(n462), .Z(n5469) );
  HS65_LS_NAND2X2 U11995 ( .A(n265), .B(n243), .Z(n5354) );
  HS65_LS_NAND2X2 U11996 ( .A(n307), .B(n285), .Z(n7061) );
  HS65_LS_NAND2X2 U11997 ( .A(n86), .B(n64), .Z(n6946) );
  HS65_LS_NAND2X2 U11998 ( .A(n699), .B(n681), .Z(n5239) );
  HS65_LS_NAND2X2 U11999 ( .A(n517), .B(n499), .Z(n6831) );
  HS65_LS_NAND2X2 U12000 ( .A(n380), .B(n388), .Z(n8275) );
  HS65_LS_OAI21X2 U12001 ( .A(n620), .B(n7710), .C(n600), .Z(n8153) );
  HS65_LS_OAI21X2 U12002 ( .A(n133), .B(n7748), .C(n113), .Z(n8185) );
  HS65_LS_NAND2X2 U12003 ( .A(n190), .B(n225), .Z(n2880) );
  HS65_LS_OAI21X2 U12004 ( .A(n210), .B(n221), .C(n189), .Z(n2876) );
  HS65_LS_OAI21X2 U12005 ( .A(n438), .B(n446), .C(n424), .Z(n3006) );
  HS65_LS_OAI21X2 U12006 ( .A(n219), .B(n214), .C(n195), .Z(n3128) );
  HS65_LS_OAI21X2 U12007 ( .A(n443), .B(n436), .C(n421), .Z(n3416) );
  HS65_LS_OAI21X2 U12008 ( .A(n172), .B(n165), .C(n157), .Z(n3295) );
  HS65_LS_OAI21X2 U12009 ( .A(n40), .B(n33), .C(n17), .Z(n4670) );
  HS65_LS_OAI21X2 U12010 ( .A(n566), .B(n559), .C(n543), .Z(n6263) );
  HS65_LS_OAI21X2 U12011 ( .A(n393), .B(n401), .C(n373), .Z(n8131) );
  HS65_LS_NAND2X2 U12012 ( .A(n345), .B(n337), .Z(n8606) );
  HS65_LS_OAI21X2 U12013 ( .A(n403), .B(n394), .C(n369), .Z(n7860) );
  HS65_LS_AOI12X2 U12014 ( .A(n600), .B(n624), .C(n8723), .Z(n8722) );
  HS65_LS_AOI12X2 U12015 ( .A(n113), .B(n137), .C(n8811), .Z(n8810) );
  HS65_LS_OAI21X2 U12016 ( .A(n669), .B(n665), .C(n650), .Z(n4252) );
  HS65_LS_OAI21X2 U12017 ( .A(n659), .B(n665), .C(n646), .Z(n4273) );
  HS65_LS_OAI21X2 U12018 ( .A(n667), .B(n660), .C(n645), .Z(n3354) );
  HS65_LS_OAI21X2 U12019 ( .A(n89), .B(n80), .C(n65), .Z(n6482) );
  HS65_LS_OAI21X2 U12020 ( .A(n310), .B(n301), .C(n286), .Z(n6596) );
  HS65_LS_OAI21X2 U12021 ( .A(n268), .B(n259), .C(n244), .Z(n4889) );
  HS65_LS_OAI21X2 U12022 ( .A(n487), .B(n478), .C(n463), .Z(n5003) );
  HS65_LS_OAI21X2 U12023 ( .A(n704), .B(n697), .C(n682), .Z(n4875) );
  HS65_LS_OAI21X2 U12024 ( .A(n522), .B(n515), .C(n500), .Z(n6468) );
  HS65_LS_OAI21X2 U12025 ( .A(n568), .B(n563), .C(n537), .Z(n7265) );
  HS65_LS_OAI21X2 U12026 ( .A(n42), .B(n37), .C(n11), .Z(n5673) );
  HS65_LS_NAND2X2 U12027 ( .A(n663), .B(n644), .Z(n3708) );
  HS65_LS_OAI21X2 U12028 ( .A(n91), .B(n85), .C(n70), .Z(n7455) );
  HS65_LS_OAI21X2 U12029 ( .A(n489), .B(n483), .C(n468), .Z(n5922) );
  HS65_LS_OAI21X2 U12030 ( .A(n312), .B(n306), .C(n291), .Z(n7514) );
  HS65_LS_OAI21X2 U12031 ( .A(n270), .B(n264), .C(n249), .Z(n5863) );
  HS65_LS_OAI21X2 U12032 ( .A(n706), .B(n701), .C(n676), .Z(n5703) );
  HS65_LS_OAI21X2 U12033 ( .A(n524), .B(n519), .C(n494), .Z(n7295) );
  HS65_LS_OAI21X2 U12034 ( .A(n165), .B(n175), .C(n143), .Z(n2926) );
  HS65_LS_NOR3AX2 U12035 ( .A(n8067), .B(n7774), .C(n8068), .Z(n8057) );
  HS65_LS_OAI21X2 U12036 ( .A(n358), .B(n7784), .C(n323), .Z(n8067) );
  HS65_LS_NAND2X2 U12037 ( .A(n399), .B(n371), .Z(n8247) );
  HS65_LS_AOI12X2 U12038 ( .A(n854), .B(n874), .C(n1188), .Z(n1187) );
  HS65_LS_AOI12X2 U12039 ( .A(n895), .B(n915), .C(n2316), .Z(n2315) );
  HS65_LS_AOI12X2 U12040 ( .A(n772), .B(n792), .C(n1940), .Z(n1939) );
  HS65_LS_AOI12X2 U12041 ( .A(n813), .B(n833), .C(n1564), .Z(n1563) );
  HS65_LS_OAI21X2 U12042 ( .A(n824), .B(n818), .C(n848), .Z(n1824) );
  HS65_LS_OAI21X2 U12043 ( .A(n906), .B(n900), .C(n930), .Z(n2576) );
  HS65_LS_NOR3AX2 U12044 ( .A(n6345), .B(n6346), .C(n6347), .Z(n6334) );
  HS65_LS_OAI21X2 U12045 ( .A(n87), .B(n6348), .C(n59), .Z(n6345) );
  HS65_LS_NOR3AX2 U12046 ( .A(n4791), .B(n4792), .C(n4793), .Z(n4780) );
  HS65_LS_OAI21X2 U12047 ( .A(n485), .B(n4794), .C(n457), .Z(n4791) );
  HS65_LS_NOR3AX2 U12048 ( .A(n6384), .B(n6385), .C(n6386), .Z(n6373) );
  HS65_LS_OAI21X2 U12049 ( .A(n308), .B(n6387), .C(n280), .Z(n6384) );
  HS65_LS_NOR3AX2 U12050 ( .A(n4752), .B(n4753), .C(n4754), .Z(n4741) );
  HS65_LS_OAI21X2 U12051 ( .A(n266), .B(n4755), .C(n238), .Z(n4752) );
  HS65_LS_NOR3AX2 U12052 ( .A(n4645), .B(n4646), .C(n4647), .Z(n4633) );
  HS65_LS_OAI21X2 U12053 ( .A(n707), .B(n4648), .C(n684), .Z(n4645) );
  HS65_LS_NOR3AX2 U12054 ( .A(n6238), .B(n6239), .C(n6240), .Z(n6226) );
  HS65_LS_OAI21X2 U12055 ( .A(n525), .B(n6241), .C(n502), .Z(n6238) );
  HS65_LS_OAI21X2 U12056 ( .A(n483), .B(n477), .C(n464), .Z(n5898) );
  HS65_LS_OAI21X2 U12057 ( .A(n264), .B(n258), .C(n245), .Z(n5839) );
  HS65_LS_OAI21X2 U12058 ( .A(n701), .B(n696), .C(n680), .Z(n5690) );
  HS65_LS_OAI21X2 U12059 ( .A(n306), .B(n300), .C(n287), .Z(n7490) );
  HS65_LS_OAI21X2 U12060 ( .A(n85), .B(n79), .C(n66), .Z(n7431) );
  HS65_LS_OAI21X2 U12061 ( .A(n519), .B(n514), .C(n498), .Z(n7282) );
  HS65_LS_OAI21X2 U12062 ( .A(n84), .B(n81), .C(n60), .Z(n6485) );
  HS65_LS_OAI21X2 U12063 ( .A(n305), .B(n302), .C(n281), .Z(n6599) );
  HS65_LS_OAI21X2 U12064 ( .A(n263), .B(n260), .C(n239), .Z(n4892) );
  HS65_LS_OAI21X2 U12065 ( .A(n482), .B(n479), .C(n458), .Z(n5006) );
  HS65_LS_OAI21X2 U12066 ( .A(n520), .B(n511), .C(n501), .Z(n6471) );
  HS65_LS_NAND2X2 U12067 ( .A(n218), .B(n197), .Z(n3465) );
  HS65_LS_OAI21X2 U12068 ( .A(n223), .B(n216), .C(n190), .Z(n4073) );
  HS65_LS_OAI21X2 U12069 ( .A(n445), .B(n441), .C(n426), .Z(n4311) );
  HS65_LS_OAI21X2 U12070 ( .A(n213), .B(n216), .C(n194), .Z(n4080) );
  HS65_LS_OAI21X2 U12071 ( .A(n435), .B(n441), .C(n422), .Z(n4332) );
  HS65_LS_OAI21X2 U12072 ( .A(n865), .B(n859), .C(n889), .Z(n1448) );
  HS65_LS_OAI21X2 U12073 ( .A(n783), .B(n777), .C(n807), .Z(n2200) );
  HS65_LS_OAI21X2 U12074 ( .A(n38), .B(n29), .C(n18), .Z(n4674) );
  HS65_LS_OAI21X2 U12075 ( .A(n564), .B(n555), .C(n544), .Z(n6267) );
  HS65_LS_OAI21X2 U12076 ( .A(n125), .B(n7891), .C(n112), .Z(n7889) );
  HS65_LS_OAI21X2 U12077 ( .A(n612), .B(n7852), .C(n599), .Z(n7850) );
  HS65_LS_OAI21X2 U12078 ( .A(n866), .B(n854), .C(n885), .Z(n1212) );
  HS65_LS_OAI21X2 U12079 ( .A(n907), .B(n895), .C(n926), .Z(n2340) );
  HS65_LS_OAI21X2 U12080 ( .A(n784), .B(n772), .C(n803), .Z(n1964) );
  HS65_LS_OAI21X2 U12081 ( .A(n825), .B(n813), .C(n844), .Z(n1588) );
  HS65_LS_OAI21X2 U12082 ( .A(n37), .B(n32), .C(n15), .Z(n5660) );
  HS65_LS_OAI21X2 U12083 ( .A(n563), .B(n558), .C(n541), .Z(n7252) );
  HS65_LS_AOI12X2 U12084 ( .A(n84), .B(n64), .C(n6948), .Z(n6947) );
  HS65_LS_AOI12X2 U12085 ( .A(n305), .B(n285), .C(n7063), .Z(n7062) );
  HS65_LS_AOI12X2 U12086 ( .A(n482), .B(n462), .C(n5471), .Z(n5470) );
  HS65_LS_AOI12X2 U12087 ( .A(n263), .B(n243), .C(n5356), .Z(n5355) );
  HS65_LS_AOI12X2 U12088 ( .A(n702), .B(n681), .C(n5241), .Z(n5240) );
  HS65_LS_AOI12X2 U12089 ( .A(n520), .B(n499), .C(n6833), .Z(n6832) );
  HS65_LS_OAI21X2 U12090 ( .A(n176), .B(n170), .C(n144), .Z(n4104) );
  HS65_LS_OAI21X2 U12091 ( .A(n167), .B(n170), .C(n149), .Z(n4111) );
  HS65_LS_AOI12X2 U12092 ( .A(n557), .B(n546), .C(n6666), .Z(n6665) );
  HS65_LS_AOI12X2 U12093 ( .A(n31), .B(n20), .C(n5073), .Z(n5072) );
  HS65_LS_AOI12X2 U12094 ( .A(n38), .B(n16), .C(n5105), .Z(n5104) );
  HS65_LS_AOI12X2 U12095 ( .A(n564), .B(n542), .C(n6698), .Z(n6697) );
  HS65_LS_OAI21X2 U12096 ( .A(n440), .B(n438), .C(n412), .Z(n3419) );
  HS65_LS_NOR3AX2 U12097 ( .A(n6161), .B(n6162), .C(n6163), .Z(n6149) );
  HS65_LS_OAI21X2 U12098 ( .A(n569), .B(n6164), .C(n546), .Z(n6161) );
  HS65_LS_NOR3AX2 U12099 ( .A(n4568), .B(n4569), .C(n4570), .Z(n4556) );
  HS65_LS_OAI21X2 U12100 ( .A(n43), .B(n4571), .C(n20), .Z(n4568) );
  HS65_LS_OAI21X2 U12101 ( .A(n398), .B(n403), .C(n374), .Z(n8134) );
  HS65_LS_OAI21X2 U12102 ( .A(n664), .B(n662), .C(n635), .Z(n3357) );
  HS65_LS_AOI12X2 U12103 ( .A(n633), .B(n661), .C(n3759), .Z(n3758) );
  HS65_LS_AOI12X2 U12104 ( .A(n82), .B(n59), .C(n6903), .Z(n6902) );
  HS65_LS_AOI12X2 U12105 ( .A(n261), .B(n238), .C(n5311), .Z(n5310) );
  HS65_LS_AOI12X2 U12106 ( .A(n480), .B(n457), .C(n5426), .Z(n5425) );
  HS65_LS_AOI12X2 U12107 ( .A(n303), .B(n280), .C(n7018), .Z(n7017) );
  HS65_LS_AOI12X2 U12108 ( .A(n695), .B(n684), .C(n5195), .Z(n5194) );
  HS65_LS_AOI12X2 U12109 ( .A(n513), .B(n502), .C(n6787), .Z(n6786) );
  HS65_LS_OAI21X2 U12110 ( .A(n671), .B(n3153), .C(n633), .Z(n3152) );
  HS65_LS_AOI12X2 U12111 ( .A(n322), .B(n8365), .C(n8366), .Z(n8364) );
  HS65_LS_NOR3AX2 U12112 ( .A(n3658), .B(n3659), .C(n3660), .Z(n3651) );
  HS65_LS_AOI12X2 U12113 ( .A(n158), .B(n166), .C(n3661), .Z(n3658) );
  HS65_LS_AOI12X2 U12114 ( .A(n376), .B(n404), .C(n8297), .Z(n8296) );
  HS65_LS_NAND3X2 U12115 ( .A(n8712), .B(n8713), .C(n8714), .Z(n8705) );
  HS65_LS_AOI12X2 U12116 ( .A(n593), .B(n606), .C(n7848), .Z(n8714) );
  HS65_LS_NAND3X2 U12117 ( .A(n8800), .B(n8801), .C(n8802), .Z(n8793) );
  HS65_LS_AOI12X2 U12118 ( .A(n106), .B(n119), .C(n7887), .Z(n8802) );
  HS65_LS_OAI21X2 U12119 ( .A(n222), .B(n2951), .C(n203), .Z(n2950) );
  HS65_LS_OAI21X2 U12120 ( .A(n447), .B(n3194), .C(n410), .Z(n3193) );
  HS65_LS_AOI12X2 U12121 ( .A(n203), .B(n212), .C(n3518), .Z(n3517) );
  HS65_LS_AOI12X2 U12122 ( .A(n571), .B(n551), .C(n6654), .Z(n6653) );
  HS65_LS_AOI12X2 U12123 ( .A(n45), .B(n25), .C(n5061), .Z(n5060) );
  HS65_LS_AOI12X2 U12124 ( .A(n915), .B(n909), .C(n2471), .Z(n2470) );
  HS65_LS_AOI12X2 U12125 ( .A(n833), .B(n827), .C(n1719), .Z(n1718) );
  HS65_LS_NOR3AX2 U12126 ( .A(n8618), .B(n8619), .C(n8620), .Z(n8611) );
  HS65_LS_AOI12X2 U12127 ( .A(n351), .B(n337), .C(n8621), .Z(n8618) );
  HS65_LS_AOI12X2 U12128 ( .A(n874), .B(n868), .C(n1343), .Z(n1342) );
  HS65_LS_AOI12X2 U12129 ( .A(n792), .B(n786), .C(n2095), .Z(n2094) );
  HS65_LS_AOI12X2 U12130 ( .A(n369), .B(n8123), .C(n8124), .Z(n8122) );
  HS65_LS_AOI12X2 U12131 ( .A(n410), .B(n437), .C(n3876), .Z(n3875) );
  HS65_LS_OAI21X2 U12132 ( .A(n36), .B(n48), .C(n12), .Z(n4586) );
  HS65_LS_OAI21X2 U12133 ( .A(n562), .B(n574), .C(n538), .Z(n6179) );
  HS65_LS_AOI12X2 U12134 ( .A(n217), .B(n197), .C(n3446), .Z(n3445) );
  HS65_LS_NOR4ABX2 U12135 ( .A(n5518), .B(n5654), .C(n5655), .D(n5486), .Z(
        n5648) );
  HS65_LS_NOR4ABX2 U12136 ( .A(n7110), .B(n7246), .C(n7247), .D(n7078), .Z(
        n7240) );
  HS65_LS_AOI12X2 U12137 ( .A(n814), .B(n834), .C(n1657), .Z(n1834) );
  HS65_LS_AOI12X2 U12138 ( .A(n896), .B(n916), .C(n2409), .Z(n2586) );
  HS65_LS_NOR4ABX2 U12139 ( .A(n7763), .B(n7764), .C(n7765), .D(n7766), .Z(
        n7749) );
  HS65_LS_AOI12X2 U12140 ( .A(n57), .B(n77), .C(n6066), .Z(n6891) );
  HS65_LS_AOI12X2 U12141 ( .A(n236), .B(n256), .C(n4473), .Z(n5299) );
  HS65_LS_AOI12X2 U12142 ( .A(n455), .B(n475), .C(n4519), .Z(n5414) );
  HS65_LS_AOI12X2 U12143 ( .A(n278), .B(n298), .C(n6112), .Z(n7006) );
  HS65_LS_AOI12X2 U12144 ( .A(n689), .B(n709), .C(n5183), .Z(n5182) );
  HS65_LS_AOI12X2 U12145 ( .A(n507), .B(n527), .C(n6775), .Z(n6774) );
  HS65_LS_AOI12X2 U12146 ( .A(n773), .B(n793), .C(n2033), .Z(n2210) );
  HS65_LS_AOI12X2 U12147 ( .A(n855), .B(n875), .C(n1281), .Z(n1458) );
  HS65_LS_NAND2X2 U12148 ( .A(n378), .B(n402), .Z(n8024) );
  HS65_LS_NAND2X2 U12149 ( .A(n154), .B(n180), .Z(n3554) );
  HS65_LS_AOI12X2 U12150 ( .A(n923), .B(n2375), .C(n2376), .Z(n2374) );
  HS65_LS_AOI12X2 U12151 ( .A(n841), .B(n1623), .C(n1624), .Z(n1622) );
  HS65_LS_AOI12X2 U12152 ( .A(n172), .B(n152), .C(n3572), .Z(n3571) );
  HS65_LS_NAND2X2 U12153 ( .A(n622), .B(n597), .Z(n7680) );
  HS65_LS_NAND2X2 U12154 ( .A(n135), .B(n110), .Z(n7718) );
  HS65_LS_AOI12X2 U12155 ( .A(n907), .B(n924), .C(n2418), .Z(n2417) );
  HS65_LS_AOI12X2 U12156 ( .A(n825), .B(n842), .C(n1666), .Z(n1665) );
  HS65_LS_AOI12X2 U12157 ( .A(n866), .B(n883), .C(n1290), .Z(n1289) );
  HS65_LS_AOI12X2 U12158 ( .A(n784), .B(n801), .C(n2042), .Z(n2041) );
  HS65_LS_OAI21X2 U12159 ( .A(n442), .B(n2861), .C(n412), .Z(n2859) );
  HS65_LS_OAI21X2 U12160 ( .A(n855), .B(n1141), .C(n885), .Z(n1139) );
  HS65_LS_OAI21X2 U12161 ( .A(n814), .B(n1517), .C(n844), .Z(n1515) );
  HS65_LS_OAI21X2 U12162 ( .A(n896), .B(n2269), .C(n926), .Z(n2267) );
  HS65_LS_OAI21X2 U12163 ( .A(n773), .B(n1893), .C(n803), .Z(n1891) );
  HS65_LS_NAND2X2 U12164 ( .A(n639), .B(n656), .Z(n3672) );
  HS65_LS_AOI12X2 U12165 ( .A(n440), .B(n420), .C(n3807), .Z(n3806) );
  HS65_LS_OAI21X2 U12166 ( .A(n666), .B(n2906), .C(n635), .Z(n2904) );
  HS65_LS_OAI21X2 U12167 ( .A(n215), .B(n3911), .C(n202), .Z(n4234) );
  HS65_LS_NAND2X2 U12168 ( .A(n160), .B(n182), .Z(n3628) );
  HS65_LS_AOI12X2 U12169 ( .A(n664), .B(n644), .C(n3690), .Z(n3689) );
  HS65_LS_NOR3AX2 U12170 ( .A(n8381), .B(n8382), .C(n8383), .Z(n8372) );
  HS65_LS_NAND2X2 U12171 ( .A(n848), .B(n819), .Z(n1682) );
  HS65_LS_NAND2X2 U12172 ( .A(n889), .B(n860), .Z(n1306) );
  HS65_LS_NAND2X2 U12173 ( .A(n930), .B(n901), .Z(n2434) );
  HS65_LS_NAND2X2 U12174 ( .A(n807), .B(n778), .Z(n2058) );
  HS65_LS_NOR3AX2 U12175 ( .A(n8025), .B(n8026), .C(n8027), .Z(n8015) );
  HS65_LS_OAI21X2 U12176 ( .A(n395), .B(n7753), .C(n376), .Z(n8025) );
  HS65_LS_OAI21X2 U12177 ( .A(n169), .B(n3921), .C(n157), .Z(n4172) );
  HS65_LS_NAND2X2 U12178 ( .A(n174), .B(n153), .Z(n3611) );
  HS65_LS_AOI12X2 U12179 ( .A(n648), .B(n3333), .C(n3334), .Z(n3332) );
  HS65_LS_NAND2X2 U12180 ( .A(n650), .B(n667), .Z(n3722) );
  HS65_LS_NAND2X2 U12181 ( .A(n394), .B(n379), .Z(n8313) );
  HS65_LS_NAND2X2 U12182 ( .A(n660), .B(n636), .Z(n3757) );
  HS65_LS_NAND2X2 U12183 ( .A(n817), .B(n840), .Z(n1717) );
  HS65_LS_NAND2X2 U12184 ( .A(n899), .B(n922), .Z(n2469) );
  HS65_LS_NAND2X2 U12185 ( .A(n356), .B(n330), .Z(n8540) );
  HS65_LS_NAND2X2 U12186 ( .A(n901), .B(n916), .Z(n2482) );
  HS65_LS_NAND2X2 U12187 ( .A(n819), .B(n834), .Z(n1730) );
  HS65_LS_NAND2X2 U12188 ( .A(n860), .B(n875), .Z(n1354) );
  HS65_LS_NAND2X2 U12189 ( .A(n778), .B(n793), .Z(n2106) );
  HS65_LS_NAND2X2 U12190 ( .A(n858), .B(n881), .Z(n1341) );
  HS65_LS_NAND2X2 U12191 ( .A(n776), .B(n799), .Z(n2093) );
  HS65_LS_NAND2X2 U12192 ( .A(n214), .B(n204), .Z(n3516) );
  HS65_LS_NAND2X2 U12193 ( .A(n394), .B(n377), .Z(n8115) );
  HS65_LS_NAND2X2 U12194 ( .A(n596), .B(n623), .Z(n8411) );
  HS65_LS_NAND2X2 U12195 ( .A(n109), .B(n136), .Z(n8471) );
  HS65_LS_NAND2X2 U12196 ( .A(n157), .B(n171), .Z(n3629) );
  HS65_LS_NAND2X2 U12197 ( .A(n670), .B(n640), .Z(n3774) );
  HS65_LS_NAND2X2 U12198 ( .A(n356), .B(n326), .Z(n8357) );
  HS65_LS_NAND2X2 U12199 ( .A(n391), .B(n377), .Z(n8294) );
  HS65_LS_NAND2X2 U12200 ( .A(n622), .B(n594), .Z(n8759) );
  HS65_LS_NAND2X2 U12201 ( .A(n135), .B(n107), .Z(n8847) );
  HS65_LS_NAND2X2 U12202 ( .A(n443), .B(n414), .Z(n3825) );
  HS65_LS_NAND2X2 U12203 ( .A(n828), .B(n843), .Z(n1750) );
  HS65_LS_NAND2X2 U12204 ( .A(n910), .B(n925), .Z(n2502) );
  HS65_LS_NAND2X2 U12205 ( .A(n869), .B(n884), .Z(n1374) );
  HS65_LS_NAND2X2 U12206 ( .A(n787), .B(n802), .Z(n2126) );
  HS65_LS_NAND2X2 U12207 ( .A(n446), .B(n416), .Z(n3891) );
  HS65_LS_NAND2X2 U12208 ( .A(n446), .B(n420), .Z(n3826) );
  HS65_LS_NAND2X2 U12209 ( .A(n221), .B(n201), .Z(n3534) );
  HS65_LS_NAND2X2 U12210 ( .A(n356), .B(n329), .Z(n8331) );
  HS65_LS_NAND2X2 U12211 ( .A(n599), .B(n615), .Z(n8697) );
  HS65_LS_NAND2X2 U12212 ( .A(n112), .B(n128), .Z(n8785) );
  HS65_LS_NAND2X2 U12213 ( .A(n899), .B(n916), .Z(n2439) );
  HS65_LS_NAND2X2 U12214 ( .A(n817), .B(n834), .Z(n1687) );
  HS65_LS_NAND2X2 U12215 ( .A(n647), .B(n659), .Z(n3732) );
  HS65_LS_NAND2X2 U12216 ( .A(n218), .B(n204), .Z(n2970) );
  HS65_LS_NAND2X2 U12217 ( .A(n213), .B(n198), .Z(n3524) );
  HS65_LS_NAND2X2 U12218 ( .A(n776), .B(n793), .Z(n2063) );
  HS65_LS_NAND2X2 U12219 ( .A(n858), .B(n875), .Z(n1311) );
  HS65_LS_AOI12X2 U12220 ( .A(n381), .B(n388), .C(n8286), .Z(n8285) );
  HS65_LS_NAND2X2 U12221 ( .A(n436), .B(n413), .Z(n3874) );
  HS65_LS_AOI12X2 U12222 ( .A(n332), .B(n348), .C(n8589), .Z(n8588) );
  HS65_LS_NAND2X2 U12223 ( .A(n660), .B(n637), .Z(n3727) );
  HS65_LS_NAND2X2 U12224 ( .A(n192), .B(n213), .Z(n3490) );
  HS65_LS_NAND2X2 U12225 ( .A(n479), .B(n456), .Z(n4991) );
  HS65_LS_NAND2X2 U12226 ( .A(n260), .B(n237), .Z(n4937) );
  HS65_LS_NAND2X2 U12227 ( .A(n302), .B(n279), .Z(n6584) );
  HS65_LS_NAND2X2 U12228 ( .A(n693), .B(n690), .Z(n4863) );
  HS65_LS_NAND2X2 U12229 ( .A(n511), .B(n508), .Z(n6456) );
  HS65_LS_NAND2X2 U12230 ( .A(n81), .B(n58), .Z(n6530) );
  HS65_LS_OAI21X2 U12231 ( .A(n461), .B(n466), .C(n480), .Z(n4522) );
  HS65_LS_OAI21X2 U12232 ( .A(n242), .B(n247), .C(n261), .Z(n4476) );
  HS65_LS_OAI21X2 U12233 ( .A(n284), .B(n289), .C(n303), .Z(n6115) );
  HS65_LS_OAI21X2 U12234 ( .A(n679), .B(n675), .C(n695), .Z(n5828) );
  HS65_LS_OAI21X2 U12235 ( .A(n497), .B(n493), .C(n513), .Z(n7420) );
  HS65_LS_OAI21X2 U12236 ( .A(n63), .B(n68), .C(n82), .Z(n6069) );
  HS65_LS_OAI21X2 U12237 ( .A(n419), .B(n424), .C(n437), .Z(n2860) );
  HS65_LS_NAND2X2 U12238 ( .A(n401), .B(n377), .Z(n8295) );
  HS65_LS_NAND2X2 U12239 ( .A(n214), .B(n198), .Z(n3485) );
  HS65_LS_NAND2X2 U12240 ( .A(n436), .B(n414), .Z(n3844) );
  HS65_LS_OAI21X2 U12241 ( .A(n14), .B(n10), .C(n31), .Z(n5766) );
  HS65_LS_OAI21X2 U12242 ( .A(n540), .B(n536), .C(n557), .Z(n7358) );
  HS65_LS_NAND2X2 U12243 ( .A(n618), .B(n601), .Z(n7647) );
  HS65_LS_NAND2X2 U12244 ( .A(n131), .B(n114), .Z(n7675) );
  HS65_LS_NAND2X2 U12245 ( .A(n29), .B(n26), .Z(n4723) );
  HS65_LS_NAND2X2 U12246 ( .A(n555), .B(n552), .Z(n6316) );
  HS65_LS_NAND2X2 U12247 ( .A(n356), .B(n318), .Z(n8362) );
  HS65_LS_NAND2X2 U12248 ( .A(n374), .B(n387), .Z(n8253) );
  HS65_LS_NAND2X2 U12249 ( .A(n412), .B(n432), .Z(n3830) );
  HS65_LS_NAND2X2 U12250 ( .A(n324), .B(n347), .Z(n8557) );
  HS65_LS_NAND2X2 U12251 ( .A(n344), .B(n326), .Z(n8599) );
  HS65_LS_NAND2X2 U12252 ( .A(n324), .B(n352), .Z(n8563) );
  HS65_LS_NAND2X2 U12253 ( .A(n32), .B(n23), .Z(n5078) );
  HS65_LS_NAND2X2 U12254 ( .A(n558), .B(n549), .Z(n6671) );
  HS65_LS_OAI21X2 U12255 ( .A(n353), .B(n343), .C(n334), .Z(n8878) );
  HS65_LS_NAND2X2 U12256 ( .A(n192), .B(n226), .Z(n3096) );
  HS65_LS_NAND2X2 U12257 ( .A(n202), .B(n226), .Z(n3471) );
  HS65_LS_OAI21X2 U12258 ( .A(n396), .B(n402), .C(n372), .Z(n8504) );
  HS65_LS_NAND2X2 U12259 ( .A(n150), .B(n166), .Z(n3259) );
  HS65_LS_NAND2X2 U12260 ( .A(n150), .B(n171), .Z(n3273) );
  HS65_LS_NAND2X2 U12261 ( .A(n439), .B(n413), .Z(n3213) );
  HS65_LS_NOR4ABX2 U12262 ( .A(n3979), .B(n3980), .C(n3981), .D(n3982), .Z(
        n3975) );
  HS65_LS_MX41X4 U12263 ( .D0(n446), .S0(n419), .D1(n413), .S1(n441), .D2(n438), .S2(n417), .D3(n415), .S3(n430), .Z(n3982) );
  HS65_LS_NOR4ABX2 U12264 ( .A(n3958), .B(n3959), .C(n3960), .D(n3961), .Z(
        n3954) );
  HS65_LS_MX41X4 U12265 ( .D0(n670), .S0(n643), .D1(n636), .S1(n665), .D2(n662), .S2(n641), .D3(n639), .S3(n654), .Z(n3961) );
  HS65_LS_NAND2X2 U12266 ( .A(n20), .B(n41), .Z(n5053) );
  HS65_LS_NAND2X2 U12267 ( .A(n546), .B(n567), .Z(n6646) );
  HS65_LS_OAI21X2 U12268 ( .A(n838), .B(n841), .C(n827), .Z(n1516) );
  HS65_LS_OAI21X2 U12269 ( .A(n920), .B(n923), .C(n909), .Z(n2268) );
  HS65_LS_NAND2X2 U12270 ( .A(n477), .B(n453), .Z(n5432) );
  HS65_LS_NAND2X2 U12271 ( .A(n258), .B(n234), .Z(n5317) );
  HS65_LS_NAND2X2 U12272 ( .A(n696), .B(n687), .Z(n5201) );
  HS65_LS_NAND2X2 U12273 ( .A(n300), .B(n276), .Z(n7024) );
  HS65_LS_NAND2X2 U12274 ( .A(n514), .B(n505), .Z(n6793) );
  HS65_LS_NAND2X2 U12275 ( .A(n79), .B(n55), .Z(n6909) );
  HS65_LS_OAI21X2 U12276 ( .A(n879), .B(n882), .C(n868), .Z(n1140) );
  HS65_LS_OAI21X2 U12277 ( .A(n797), .B(n800), .C(n786), .Z(n1892) );
  HS65_LS_NAND2X2 U12278 ( .A(n65), .B(n91), .Z(n6886) );
  HS65_LS_NAND2X2 U12279 ( .A(n463), .B(n489), .Z(n5409) );
  HS65_LS_NAND2X2 U12280 ( .A(n286), .B(n312), .Z(n7001) );
  HS65_LS_NAND2X2 U12281 ( .A(n244), .B(n270), .Z(n5294) );
  HS65_LS_NAND2X2 U12282 ( .A(n682), .B(n706), .Z(n5177) );
  HS65_LS_NAND2X2 U12283 ( .A(n500), .B(n524), .Z(n6769) );
  HS65_LS_NAND2X2 U12284 ( .A(n599), .B(n616), .Z(n8727) );
  HS65_LS_NAND2X2 U12285 ( .A(n112), .B(n129), .Z(n8815) );
  HS65_LS_OAI21X2 U12286 ( .A(n335), .B(n322), .C(n345), .Z(n8643) );
  HS65_LS_OAI21X2 U12287 ( .A(n370), .B(n369), .C(n404), .Z(n8675) );
  HS65_LS_NAND2X2 U12288 ( .A(n423), .B(n432), .Z(n3387) );
  HS65_LS_OAI21X2 U12289 ( .A(n586), .B(n585), .C(n606), .Z(n7805) );
  HS65_LS_OAI21X2 U12290 ( .A(n99), .B(n98), .C(n119), .Z(n7905) );
  HS65_LS_NAND2X2 U12291 ( .A(n380), .B(n399), .Z(n8317) );
  HS65_LS_NAND2X2 U12292 ( .A(n615), .B(n585), .Z(n7704) );
  HS65_LS_NAND2X2 U12293 ( .A(n128), .B(n98), .Z(n7742) );
  HS65_LS_OAI21X2 U12294 ( .A(n643), .B(n648), .C(n661), .Z(n2905) );
  HS65_LS_NAND2X2 U12295 ( .A(n659), .B(n637), .Z(n3765) );
  HS65_LS_OAI21X2 U12296 ( .A(n150), .B(n148), .C(n179), .Z(n4133) );
  HS65_LS_OAI21X2 U12297 ( .A(n373), .B(n370), .C(n388), .Z(n8970) );
  HS65_LS_NAND3X2 U12298 ( .A(n4723), .B(n4724), .C(n4725), .Z(n4707) );
  HS65_LS_AOI12X2 U12299 ( .A(n10), .B(n4726), .C(n4727), .Z(n4725) );
  HS65_LS_NAND3X2 U12300 ( .A(n6316), .B(n6317), .C(n6318), .Z(n6300) );
  HS65_LS_AOI12X2 U12301 ( .A(n536), .B(n6319), .C(n6320), .Z(n6318) );
  HS65_LS_OAI21X2 U12302 ( .A(n336), .B(n335), .C(n348), .Z(n8910) );
  HS65_LS_OAI21X2 U12303 ( .A(n11), .B(n10), .C(n42), .Z(n4585) );
  HS65_LS_OAI21X2 U12304 ( .A(n537), .B(n536), .C(n568), .Z(n6178) );
  HS65_LS_OAI21X2 U12305 ( .A(n468), .B(n466), .C(n489), .Z(n4808) );
  HS65_LS_AOI12X2 U12306 ( .A(n155), .B(n179), .C(n3645), .Z(n3644) );
  HS65_LS_OAI21X2 U12307 ( .A(n929), .B(n923), .C(n903), .Z(n2392) );
  HS65_LS_OAI21X2 U12308 ( .A(n847), .B(n841), .C(n821), .Z(n1640) );
  HS65_LS_NAND2X2 U12309 ( .A(n374), .B(n393), .Z(n8299) );
  HS65_LS_NOR4ABX2 U12310 ( .A(n8726), .B(n8727), .C(n7836), .D(n8728), .Z(
        n8717) );
  HS65_LS_NOR4ABX2 U12311 ( .A(n8814), .B(n8815), .C(n7935), .D(n8816), .Z(
        n8805) );
  HS65_LS_OAI21X2 U12312 ( .A(n888), .B(n882), .C(n862), .Z(n1264) );
  HS65_LS_OAI21X2 U12313 ( .A(n806), .B(n800), .C(n780), .Z(n2016) );
  HS65_LS_NAND2X2 U12314 ( .A(n104), .B(n126), .Z(n8828) );
  HS65_LS_NAND2X2 U12315 ( .A(n591), .B(n613), .Z(n8740) );
  HS65_LS_OAI21X2 U12316 ( .A(n327), .B(n322), .C(n352), .Z(n8380) );
  HS65_LS_NOR4ABX2 U12317 ( .A(n7806), .B(n7807), .C(n7808), .D(n7809), .Z(
        n7795) );
  HS65_LS_NOR4ABX2 U12318 ( .A(n7906), .B(n7907), .C(n7908), .D(n7909), .Z(
        n7895) );
  HS65_LS_OAI21X2 U12319 ( .A(n634), .B(n648), .C(n663), .Z(n3350) );
  HS65_LS_NAND2X2 U12320 ( .A(n857), .B(n888), .Z(n1179) );
  HS65_LS_NAND2X2 U12321 ( .A(n775), .B(n806), .Z(n1931) );
  HS65_LS_NAND2X2 U12322 ( .A(n898), .B(n929), .Z(n2307) );
  HS65_LS_NAND2X2 U12323 ( .A(n816), .B(n847), .Z(n1555) );
  HS65_LS_OAI21X2 U12324 ( .A(n650), .B(n648), .C(n669), .Z(n3171) );
  HS65_LS_NAND2X2 U12325 ( .A(n217), .B(n191), .Z(n3097) );
  HS65_LS_NOR4ABX2 U12326 ( .A(n6905), .B(n6914), .C(n6883), .D(n6522), .Z(
        n7469) );
  HS65_LS_NOR4ABX2 U12327 ( .A(n5428), .B(n5437), .C(n5406), .D(n4983), .Z(
        n5936) );
  HS65_LS_NOR4ABX2 U12328 ( .A(n7020), .B(n7029), .C(n6998), .D(n6576), .Z(
        n7528) );
  HS65_LS_NOR4ABX2 U12329 ( .A(n5313), .B(n5322), .C(n5291), .D(n4929), .Z(
        n5877) );
  HS65_LS_NOR4ABX2 U12330 ( .A(n5197), .B(n5206), .C(n5174), .D(n4853), .Z(
        n5773) );
  HS65_LS_NOR4ABX2 U12331 ( .A(n6789), .B(n6798), .C(n6766), .D(n6446), .Z(
        n7365) );
  HS65_LS_NAND2X2 U12332 ( .A(n346), .B(n322), .Z(n8587) );
  HS65_LS_NOR4ABX2 U12333 ( .A(n6667), .B(n6678), .C(n6645), .D(n6306), .Z(
        n7303) );
  HS65_LS_NOR4ABX2 U12334 ( .A(n5074), .B(n5085), .C(n5052), .D(n4713), .Z(
        n5711) );
  HS65_LS_NAND2X2 U12335 ( .A(n147), .B(n179), .Z(n3634) );
  HS65_LS_NOR4ABX2 U12336 ( .A(n4074), .B(n4060), .C(n3935), .D(n4201), .Z(
        n4197) );
  HS65_LS_MX41X4 U12337 ( .D0(n221), .S0(n193), .D1(n204), .S1(n216), .D2(n210), .S2(n200), .D3(n199), .S3(n227), .Z(n4201) );
  HS65_LS_NOR4ABX2 U12338 ( .A(n5457), .B(n4991), .C(n5380), .D(n4792), .Z(
        n5635) );
  HS65_LS_NOR4ABX2 U12339 ( .A(n5342), .B(n4937), .C(n5265), .D(n4753), .Z(
        n5608) );
  HS65_LS_NOR4ABX2 U12340 ( .A(n7049), .B(n6584), .C(n6972), .D(n6385), .Z(
        n7227) );
  HS65_LS_NOR4ABX2 U12341 ( .A(n5226), .B(n4863), .C(n5147), .D(n4646), .Z(
        n5801) );
  HS65_LS_NOR4ABX2 U12342 ( .A(n6818), .B(n6456), .C(n6739), .D(n6239), .Z(
        n7393) );
  HS65_LS_NOR4ABX2 U12343 ( .A(n6934), .B(n6530), .C(n6857), .D(n6346), .Z(
        n7200) );
  HS65_LS_NOR4ABX2 U12344 ( .A(n3523), .B(n3465), .C(n3504), .D(n3099), .Z(
        n4180) );
  HS65_LSS_XOR2X3 U12345 ( .A(n2639), .B(n2728), .Z(n2704) );
  HS65_LS_NOR4ABX2 U12346 ( .A(n3891), .B(n3825), .C(n3197), .D(n3385), .Z(
        n4043) );
  HS65_LS_NOR4ABX2 U12347 ( .A(n3523), .B(n3524), .C(n3525), .D(n3526), .Z(
        n3511) );
  HS65_LS_NAND4ABX3 U12348 ( .A(n3356), .B(n3673), .C(n3172), .D(n3747), .Z(
        n4261) );
  HS65_LS_NAND2X2 U12349 ( .A(n606), .B(n592), .Z(n7976) );
  HS65_LS_NAND2X2 U12350 ( .A(n119), .B(n105), .Z(n7989) );
  HS65_LS_NOR4ABX2 U12351 ( .A(n3774), .B(n3155), .C(n3707), .D(n3323), .Z(
        n4019) );
  HS65_LS_NAND2X2 U12352 ( .A(n375), .B(n397), .Z(n8112) );
  HS65_LS_NAND2X2 U12353 ( .A(n411), .B(n442), .Z(n3384) );
  HS65_LS_OAI21X2 U12354 ( .A(n484), .B(n485), .C(n457), .Z(n5567) );
  HS65_LS_OAI21X2 U12355 ( .A(n265), .B(n266), .C(n238), .Z(n5546) );
  HS65_LS_OAI21X2 U12356 ( .A(n307), .B(n308), .C(n280), .Z(n7159) );
  HS65_LS_OAI21X2 U12357 ( .A(n699), .B(n707), .C(n684), .Z(n5821) );
  HS65_LS_OAI21X2 U12358 ( .A(n517), .B(n525), .C(n502), .Z(n7413) );
  HS65_LS_OAI21X2 U12359 ( .A(n86), .B(n87), .C(n59), .Z(n7138) );
  HS65_LS_OAI21X2 U12360 ( .A(n397), .B(n395), .C(n376), .Z(n8665) );
  HS65_LS_OAI21X2 U12361 ( .A(n929), .B(n922), .C(n901), .Z(n2302) );
  HS65_LS_OAI21X2 U12362 ( .A(n847), .B(n840), .C(n819), .Z(n1550) );
  HS65_LS_OAI21X2 U12363 ( .A(n614), .B(n625), .C(n584), .Z(n9049) );
  HS65_LS_OAI21X2 U12364 ( .A(n127), .B(n138), .C(n97), .Z(n9107) );
  HS65_LS_OAI21X2 U12365 ( .A(n616), .B(n614), .C(n583), .Z(n7643) );
  HS65_LS_OAI21X2 U12366 ( .A(n129), .B(n127), .C(n96), .Z(n7671) );
  HS65_LS_NAND2X2 U12367 ( .A(n109), .B(n126), .Z(n7924) );
  HS65_LS_NAND2X2 U12368 ( .A(n596), .B(n613), .Z(n7825) );
  HS65_LS_NAND2X2 U12369 ( .A(n583), .B(n625), .Z(n8712) );
  HS65_LS_NAND2X2 U12370 ( .A(n96), .B(n138), .Z(n8800) );
  HS65_LS_NAND2X2 U12371 ( .A(n634), .B(n666), .Z(n3322) );
  HS65_LS_NAND2X2 U12372 ( .A(n205), .B(n215), .Z(n3093) );
  HS65_LS_OAI21X2 U12373 ( .A(n888), .B(n881), .C(n860), .Z(n1174) );
  HS65_LS_OAI21X2 U12374 ( .A(n806), .B(n799), .C(n778), .Z(n1926) );
  HS65_LS_NOR4ABX2 U12375 ( .A(n8298), .B(n8299), .C(n8300), .D(n8301), .Z(
        n8291) );
  HS65_LS_OAI21X2 U12376 ( .A(n442), .B(n447), .C(n410), .Z(n3978) );
  HS65_LS_NOR4ABX2 U12377 ( .A(n2970), .B(n3506), .C(n3130), .D(n3429), .Z(
        n4217) );
  HS65_LS_NAND2X2 U12378 ( .A(n806), .B(n773), .Z(n1988) );
  HS65_LS_NAND2X2 U12379 ( .A(n888), .B(n855), .Z(n1236) );
  HS65_LS_NAND2X2 U12380 ( .A(n847), .B(n814), .Z(n1612) );
  HS65_LS_NAND2X2 U12381 ( .A(n929), .B(n896), .Z(n2364) );
  HS65_LS_OAI21X2 U12382 ( .A(n666), .B(n671), .C(n633), .Z(n3957) );
  HS65_LS_NAND2X2 U12383 ( .A(n460), .B(n472), .Z(n5394) );
  HS65_LS_NAND2X2 U12384 ( .A(n241), .B(n253), .Z(n5279) );
  HS65_LS_NAND2X2 U12385 ( .A(n283), .B(n295), .Z(n6986) );
  HS65_LS_NAND2X2 U12386 ( .A(n686), .B(n712), .Z(n5162) );
  HS65_LS_NAND2X2 U12387 ( .A(n504), .B(n530), .Z(n6754) );
  HS65_LS_NAND2X2 U12388 ( .A(n62), .B(n74), .Z(n6871) );
  HS65_LS_NOR4ABX2 U12389 ( .A(n3283), .B(n3648), .C(n3040), .D(n3257), .Z(
        n4151) );
  HS65_LS_NAND2X2 U12390 ( .A(n147), .B(n182), .Z(n3635) );
  HS65_LS_NOR4ABX2 U12391 ( .A(n5120), .B(n4723), .C(n5025), .D(n4569), .Z(
        n5739) );
  HS65_LS_NOR4ABX2 U12392 ( .A(n6713), .B(n6316), .C(n6618), .D(n6162), .Z(
        n7331) );
  HS65_LS_NAND2X2 U12393 ( .A(n929), .B(n908), .Z(n2443) );
  HS65_LS_NAND2X2 U12394 ( .A(n847), .B(n826), .Z(n1691) );
  HS65_LS_NAND2X2 U12395 ( .A(n334), .B(n352), .Z(n8583) );
  HS65_LS_NOR4ABX2 U12396 ( .A(n3764), .B(n3765), .C(n3766), .D(n3767), .Z(
        n3752) );
  HS65_LS_NAND2X2 U12397 ( .A(n888), .B(n867), .Z(n1315) );
  HS65_LS_NAND2X2 U12398 ( .A(n223), .B(n204), .Z(n3515) );
  HS65_LS_NAND2X2 U12399 ( .A(n669), .B(n636), .Z(n3756) );
  HS65_LS_NOR4ABX2 U12400 ( .A(n2107), .B(n1912), .C(n2056), .D(n2124), .Z(
        n2206) );
  HS65_LS_NOR4ABX2 U12401 ( .A(n1355), .B(n1160), .C(n1304), .D(n1372), .Z(
        n1454) );
  HS65_LS_NOR4ABX2 U12402 ( .A(n1731), .B(n1536), .C(n1680), .D(n1748), .Z(
        n1830) );
  HS65_LS_NOR4ABX2 U12403 ( .A(n2483), .B(n2288), .C(n2432), .D(n2500), .Z(
        n2582) );
  HS65_LS_NAND2X2 U12404 ( .A(n109), .B(n132), .Z(n8834) );
  HS65_LS_NAND2X2 U12405 ( .A(n596), .B(n619), .Z(n8746) );
  HS65_LS_NAND2X2 U12406 ( .A(n155), .B(n181), .Z(n3565) );
  HS65_LS_NOR4ABX2 U12407 ( .A(n8606), .B(n8607), .C(n8608), .D(n8609), .Z(
        n8594) );
  HS65_LS_NAND2X2 U12408 ( .A(n598), .B(n609), .Z(n8701) );
  HS65_LS_NAND2X2 U12409 ( .A(n111), .B(n122), .Z(n8789) );
  HS65_LS_NAND2X2 U12410 ( .A(n806), .B(n785), .Z(n2067) );
  HS65_LS_NAND3AX3 U12411 ( .A(n2303), .B(n2304), .C(n2305), .Z(n2297) );
  HS65_LS_OAI21X2 U12412 ( .A(n897), .B(n2306), .C(n915), .Z(n2305) );
  HS65_LS_NAND3AX3 U12413 ( .A(n1551), .B(n1552), .C(n1553), .Z(n1545) );
  HS65_LS_OAI21X2 U12414 ( .A(n815), .B(n1554), .C(n833), .Z(n1553) );
  HS65_LS_NAND3AX3 U12415 ( .A(n1175), .B(n1176), .C(n1177), .Z(n1169) );
  HS65_LS_OAI21X2 U12416 ( .A(n856), .B(n1178), .C(n874), .Z(n1177) );
  HS65_LS_NAND3AX3 U12417 ( .A(n1927), .B(n1928), .C(n1929), .Z(n1921) );
  HS65_LS_OAI21X2 U12418 ( .A(n774), .B(n1930), .C(n792), .Z(n1929) );
  HS65_LS_NOR4ABX2 U12419 ( .A(n3104), .B(n3515), .C(n3488), .D(n3508), .Z(
        n4077) );
  HS65_LS_NAND2X2 U12420 ( .A(n62), .B(n80), .Z(n6904) );
  HS65_LS_NAND2X2 U12421 ( .A(n241), .B(n259), .Z(n5312) );
  HS65_LS_NAND2X2 U12422 ( .A(n460), .B(n478), .Z(n5427) );
  HS65_LS_NAND2X2 U12423 ( .A(n283), .B(n301), .Z(n7019) );
  HS65_LS_NAND2X2 U12424 ( .A(n686), .B(n697), .Z(n5196) );
  HS65_LS_NAND2X2 U12425 ( .A(n504), .B(n515), .Z(n6788) );
  HS65_LS_NOR4ABX2 U12426 ( .A(n6908), .B(n6909), .C(n6910), .D(n6911), .Z(
        n6896) );
  HS65_LS_NOR4ABX2 U12427 ( .A(n5316), .B(n5317), .C(n5318), .D(n5319), .Z(
        n5304) );
  HS65_LS_NOR4ABX2 U12428 ( .A(n5431), .B(n5432), .C(n5433), .D(n5434), .Z(
        n5419) );
  HS65_LS_NOR4ABX2 U12429 ( .A(n7023), .B(n7024), .C(n7025), .D(n7026), .Z(
        n7011) );
  HS65_LS_NOR4ABX2 U12430 ( .A(n5200), .B(n5201), .C(n5202), .D(n5203), .Z(
        n5188) );
  HS65_LS_NOR4ABX2 U12431 ( .A(n6792), .B(n6793), .C(n6794), .D(n6795), .Z(
        n6780) );
  HS65_LS_OAI21X2 U12432 ( .A(n98), .B(n104), .C(n137), .Z(n7890) );
  HS65_LS_OAI21X2 U12433 ( .A(n585), .B(n591), .C(n624), .Z(n7851) );
  HS65_LS_NAND2X2 U12434 ( .A(n347), .B(n330), .Z(n8370) );
  HS65_LS_OAI21X2 U12435 ( .A(n205), .B(n204), .C(n219), .Z(n2947) );
  HS65_LS_OAI21X2 U12436 ( .A(n634), .B(n636), .C(n667), .Z(n3149) );
  HS65_LS_NAND2X2 U12437 ( .A(n619), .B(n598), .Z(n7698) );
  HS65_LS_NAND2X2 U12438 ( .A(n132), .B(n111), .Z(n7736) );
  HS65_LS_NOR4ABX2 U12439 ( .A(n4149), .B(n3583), .C(n3568), .D(n3593), .Z(
        n4144) );
  HS65_LS_OAI21X2 U12440 ( .A(n149), .B(n147), .C(n166), .Z(n4149) );
  HS65_LS_NAND2X2 U12441 ( .A(n564), .B(n541), .Z(n6643) );
  HS65_LS_NAND2X2 U12442 ( .A(n38), .B(n15), .Z(n5050) );
  HS65_LS_NOR4ABX2 U12443 ( .A(n3617), .B(n3296), .C(n3664), .D(n3646), .Z(
        n3999) );
  HS65_LS_NAND4ABX3 U12444 ( .A(n8133), .B(n8210), .C(n8008), .D(n8280), .Z(
        n8959) );
  HS65_LS_NAND2X2 U12445 ( .A(n357), .B(n331), .Z(n8551) );
  HS65_LS_OAI21X2 U12446 ( .A(n411), .B(n413), .C(n443), .Z(n3190) );
  HS65_LS_NOR4ABX2 U12447 ( .A(n8369), .B(n8381), .C(n8582), .D(n8615), .Z(
        n8923) );
  HS65_LS_NAND2X2 U12448 ( .A(n370), .B(n402), .Z(n8266) );
  HS65_LS_NOR4ABX2 U12449 ( .A(n8313), .B(n8024), .C(n8113), .D(n8246), .Z(
        n8990) );
  HS65_LS_NAND2X2 U12450 ( .A(n455), .B(n481), .Z(n5431) );
  HS65_LS_NAND2X2 U12451 ( .A(n236), .B(n262), .Z(n5316) );
  HS65_LS_NAND2X2 U12452 ( .A(n278), .B(n304), .Z(n7023) );
  HS65_LS_NAND2X2 U12453 ( .A(n689), .B(n700), .Z(n5200) );
  HS65_LS_NAND2X2 U12454 ( .A(n57), .B(n83), .Z(n6908) );
  HS65_LS_NAND2X2 U12455 ( .A(n507), .B(n518), .Z(n6792) );
  HS65_LS_OAI21X2 U12456 ( .A(n375), .B(n377), .C(n393), .Z(n8020) );
  HS65_LS_OAI21X2 U12457 ( .A(n327), .B(n326), .C(n357), .Z(n8062) );
  HS65_LS_NOR4ABX2 U12458 ( .A(n8362), .B(n8331), .C(n8572), .D(n8590), .Z(
        n8931) );
  HS65_LS_NOR4ABX2 U12459 ( .A(n3213), .B(n3864), .C(n3418), .D(n3790), .Z(
        n4320) );
  HS65_LS_NAND2X2 U12460 ( .A(n664), .B(n640), .Z(n3683) );
  HS65_LS_NAND2X2 U12461 ( .A(n591), .B(n609), .Z(n8716) );
  HS65_LS_NAND2X2 U12462 ( .A(n104), .B(n122), .Z(n8804) );
  HS65_LS_NAND2X2 U12463 ( .A(n548), .B(n559), .Z(n6668) );
  HS65_LS_NAND2X2 U12464 ( .A(n22), .B(n33), .Z(n5075) );
  HS65_LS_NAND2X2 U12465 ( .A(n828), .B(n844), .Z(n1724) );
  HS65_LS_NAND2X2 U12466 ( .A(n910), .B(n926), .Z(n2476) );
  HS65_LS_NAND2X2 U12467 ( .A(n387), .B(n379), .Z(n8128) );
  HS65_LS_NAND2X2 U12468 ( .A(n598), .B(n618), .Z(n8726) );
  HS65_LS_NAND2X2 U12469 ( .A(n111), .B(n131), .Z(n8814) );
  HS65_LS_OAI21X2 U12470 ( .A(n601), .B(n598), .C(n616), .Z(n8151) );
  HS65_LS_OAI21X2 U12471 ( .A(n114), .B(n111), .C(n129), .Z(n8183) );
  HS65_LS_NAND2X2 U12472 ( .A(n869), .B(n885), .Z(n1348) );
  HS65_LS_NAND2X2 U12473 ( .A(n787), .B(n803), .Z(n2100) );
  HS65_LS_NAND2X2 U12474 ( .A(n148), .B(n167), .Z(n3617) );
  HS65_LS_NAND2X2 U12475 ( .A(n374), .B(n394), .Z(n8303) );
  HS65_LS_NAND2X2 U12476 ( .A(n373), .B(n396), .Z(n8234) );
  HS65_LS_NOR4ABX2 U12477 ( .A(n8155), .B(n7800), .C(n7708), .D(n8156), .Z(
        n8146) );
  HS65_LS_NOR4ABX2 U12478 ( .A(n8187), .B(n7900), .C(n7746), .D(n8188), .Z(
        n8178) );
  HS65_LS_NOR4ABX2 U12479 ( .A(n6949), .B(n6950), .C(n6951), .D(n6952), .Z(
        n6942) );
  HS65_LS_NOR4ABX2 U12480 ( .A(n7064), .B(n7065), .C(n7066), .D(n7067), .Z(
        n7057) );
  HS65_LS_NOR4ABX2 U12481 ( .A(n5472), .B(n5473), .C(n5474), .D(n5475), .Z(
        n5465) );
  HS65_LS_NOR4ABX2 U12482 ( .A(n5357), .B(n5358), .C(n5359), .D(n5360), .Z(
        n5350) );
  HS65_LS_NOR4ABX2 U12483 ( .A(n5242), .B(n5243), .C(n5244), .D(n5245), .Z(
        n5235) );
  HS65_LS_NOR4ABX2 U12484 ( .A(n6834), .B(n6835), .C(n6836), .D(n6837), .Z(
        n6827) );
  HS65_LS_NAND2X2 U12485 ( .A(n446), .B(n412), .Z(n3881) );
  HS65_LS_NAND2X2 U12486 ( .A(n324), .B(n356), .Z(n8607) );
  HS65_LS_NAND2X2 U12487 ( .A(n866), .B(n884), .Z(n1283) );
  HS65_LS_NAND2X2 U12488 ( .A(n784), .B(n802), .Z(n2035) );
  HS65_LS_NAND2X2 U12489 ( .A(n907), .B(n925), .Z(n2411) );
  HS65_LS_NAND2X2 U12490 ( .A(n825), .B(n843), .Z(n1659) );
  HS65_LS_OAI21X2 U12491 ( .A(n61), .B(n62), .C(n89), .Z(n6340) );
  HS65_LS_OAI21X2 U12492 ( .A(n459), .B(n460), .C(n487), .Z(n4786) );
  HS65_LS_OAI21X2 U12493 ( .A(n282), .B(n283), .C(n310), .Z(n6379) );
  HS65_LS_OAI21X2 U12494 ( .A(n240), .B(n241), .C(n268), .Z(n4747) );
  HS65_LS_OAI21X2 U12495 ( .A(n685), .B(n686), .C(n704), .Z(n4640) );
  HS65_LS_OAI21X2 U12496 ( .A(n503), .B(n504), .C(n522), .Z(n6233) );
  HS65_LS_NOR4ABX2 U12497 ( .A(n8303), .B(n8247), .C(n8282), .D(n8118), .Z(
        n8967) );
  HS65_LS_NOR4ABX2 U12498 ( .A(n2952), .B(n2953), .C(n2954), .D(n2955), .Z(
        n2940) );
  HS65_LS_NAND4ABX3 U12499 ( .A(n8329), .B(n8516), .C(n8050), .D(n8584), .Z(
        n8899) );
  HS65_LS_NAND2X2 U12500 ( .A(n351), .B(n330), .Z(n8622) );
  HS65_LS_NAND2X2 U12501 ( .A(n411), .B(n431), .Z(n3848) );
  HS65_LS_OAI21X2 U12502 ( .A(n25), .B(n4693), .C(n29), .Z(n4702) );
  HS65_LS_OAI21X2 U12503 ( .A(n551), .B(n6286), .C(n555), .Z(n6295) );
  HS65_LS_NAND2X2 U12504 ( .A(n670), .B(n635), .Z(n3764) );
  HS65_LS_NOR4ABX2 U12505 ( .A(n3731), .B(n3358), .C(n3759), .D(n3742), .Z(
        n4024) );
  HS65_LS_NAND2X2 U12506 ( .A(n221), .B(n202), .Z(n3523) );
  HS65_LS_OAI21X2 U12507 ( .A(n57), .B(n6503), .C(n81), .Z(n6511) );
  HS65_LS_OAI21X2 U12508 ( .A(n278), .B(n6557), .C(n302), .Z(n6565) );
  HS65_LS_OAI21X2 U12509 ( .A(n455), .B(n4964), .C(n479), .Z(n4972) );
  HS65_LS_OAI21X2 U12510 ( .A(n236), .B(n4910), .C(n260), .Z(n4918) );
  HS65_LS_OAI21X2 U12511 ( .A(n689), .B(n4833), .C(n693), .Z(n4842) );
  HS65_LS_OAI21X2 U12512 ( .A(n507), .B(n6426), .C(n511), .Z(n6435) );
  HS65_LS_NAND2X2 U12513 ( .A(n423), .B(n430), .Z(n3196) );
  HS65_LS_NOR4ABX2 U12514 ( .A(n2476), .B(n2477), .C(n2478), .D(n2479), .Z(
        n2464) );
  HS65_LS_NOR4ABX2 U12515 ( .A(n1724), .B(n1725), .C(n1726), .D(n1727), .Z(
        n1712) );
  HS65_LS_NAND2X2 U12516 ( .A(n639), .B(n659), .Z(n3155) );
  HS65_LS_NAND2X2 U12517 ( .A(n818), .B(n846), .Z(n1656) );
  HS65_LS_NAND2X2 U12518 ( .A(n900), .B(n928), .Z(n2408) );
  HS65_LS_NOR4ABX2 U12519 ( .A(n1348), .B(n1349), .C(n1350), .D(n1351), .Z(
        n1336) );
  HS65_LS_NOR4ABX2 U12520 ( .A(n2100), .B(n2101), .C(n2102), .D(n2103), .Z(
        n2088) );
  HS65_LS_NOR4ABX2 U12521 ( .A(n3154), .B(n3155), .C(n3156), .D(n3157), .Z(
        n3143) );
  HS65_LS_NAND2X2 U12522 ( .A(n482), .B(n456), .Z(n5476) );
  HS65_LS_NAND2X2 U12523 ( .A(n263), .B(n237), .Z(n5361) );
  HS65_LS_NAND2X2 U12524 ( .A(n702), .B(n690), .Z(n5246) );
  HS65_LS_NAND2X2 U12525 ( .A(n38), .B(n26), .Z(n5110) );
  HS65_LS_NAND2X2 U12526 ( .A(n305), .B(n279), .Z(n7068) );
  HS65_LS_NAND2X2 U12527 ( .A(n520), .B(n508), .Z(n6838) );
  HS65_LS_NAND2X2 U12528 ( .A(n84), .B(n58), .Z(n6953) );
  HS65_LS_NAND2X2 U12529 ( .A(n564), .B(n552), .Z(n6703) );
  HS65_LS_NAND2X2 U12530 ( .A(n157), .B(n175), .Z(n3662) );
  HS65_LS_NAND2X2 U12531 ( .A(n777), .B(n805), .Z(n2032) );
  HS65_LS_NAND2X2 U12532 ( .A(n859), .B(n887), .Z(n1280) );
  HS65_LS_NOR4ABX2 U12533 ( .A(n6531), .B(n6486), .C(n6873), .D(n6894), .Z(
        n7206) );
  HS65_LS_NOR4ABX2 U12534 ( .A(n6457), .B(n6472), .C(n6756), .D(n6778), .Z(
        n7177) );
  HS65_LS_NOR4ABX2 U12535 ( .A(n4864), .B(n4879), .C(n5164), .D(n5186), .Z(
        n5585) );
  HS65_LS_NOR4ABX2 U12536 ( .A(n4992), .B(n5007), .C(n5396), .D(n5417), .Z(
        n5641) );
  HS65_LS_NOR4ABX2 U12537 ( .A(n6585), .B(n6600), .C(n6988), .D(n7009), .Z(
        n7233) );
  HS65_LS_NOR4ABX2 U12538 ( .A(n4938), .B(n4893), .C(n5281), .D(n5302), .Z(
        n5614) );
  HS65_LSS_XOR2X3 U12539 ( .A(n2822), .B(n2798), .Z(n5958) );
  HS65_LS_NOR4ABX2 U12540 ( .A(n1692), .B(n1589), .C(n1719), .D(n1702), .Z(
        n1801) );
  HS65_LS_NOR4ABX2 U12541 ( .A(n2444), .B(n2341), .C(n2471), .D(n2454), .Z(
        n2553) );
  HS65_LS_NAND2X2 U12542 ( .A(n199), .B(n213), .Z(n2953) );
  HS65_LS_NOR4ABX2 U12543 ( .A(n3881), .B(n3882), .C(n3883), .D(n3884), .Z(
        n3869) );
  HS65_LS_NOR4ABX2 U12544 ( .A(n5106), .B(n5107), .C(n5108), .D(n5109), .Z(
        n5099) );
  HS65_LS_NOR4ABX2 U12545 ( .A(n6699), .B(n6700), .C(n6701), .D(n6702), .Z(
        n6692) );
  HS65_LS_NAND2X2 U12546 ( .A(n440), .B(n416), .Z(n3800) );
  HS65_LS_NOR4ABX2 U12547 ( .A(n2068), .B(n1965), .C(n2095), .D(n2078), .Z(
        n2177) );
  HS65_LS_NOR4ABX2 U12548 ( .A(n1316), .B(n1213), .C(n1343), .D(n1326), .Z(
        n1425) );
  HS65_LS_NOR4ABX2 U12549 ( .A(n8607), .B(n8358), .C(n8550), .D(n8586), .Z(
        n8907) );
  HS65_LS_NOR4ABX2 U12550 ( .A(n8557), .B(n8599), .C(n8524), .D(n8592), .Z(
        n8902) );
  HS65_LS_NAND2X2 U12551 ( .A(n544), .B(n567), .Z(n6667) );
  HS65_LS_NAND2X2 U12552 ( .A(n18), .B(n41), .Z(n5074) );
  HS65_LS_NAND2X2 U12553 ( .A(n174), .B(n144), .Z(n3616) );
  HS65_LS_NAND2X2 U12554 ( .A(n182), .B(n157), .Z(n3663) );
  HS65_LS_NOR4ABX2 U12555 ( .A(n3489), .B(n3132), .C(n3518), .D(n3501), .Z(
        n3937) );
  HS65_LS_NAND2X2 U12556 ( .A(n921), .B(n903), .Z(n2473) );
  HS65_LS_NAND2X2 U12557 ( .A(n839), .B(n821), .Z(n1721) );
  HS65_LS_NAND2X2 U12558 ( .A(n441), .B(n421), .Z(n3797) );
  HS65_LS_NAND2X2 U12559 ( .A(n897), .B(n928), .Z(n2368) );
  HS65_LS_NAND2X2 U12560 ( .A(n815), .B(n846), .Z(n1616) );
  HS65_LS_NAND2X2 U12561 ( .A(n332), .B(n349), .Z(n8623) );
  HS65_LS_NAND2X2 U12562 ( .A(n880), .B(n862), .Z(n1345) );
  HS65_LS_NAND2X2 U12563 ( .A(n798), .B(n780), .Z(n2097) );
  HS65_LS_NAND2X2 U12564 ( .A(n856), .B(n887), .Z(n1240) );
  HS65_LS_NAND2X2 U12565 ( .A(n774), .B(n805), .Z(n1992) );
  HS65_LS_NAND2X2 U12566 ( .A(n665), .B(n645), .Z(n3680) );
  HS65_LS_NAND2X2 U12567 ( .A(n200), .B(n218), .Z(n3520) );
  HS65_LS_NAND2X2 U12568 ( .A(n60), .B(n88), .Z(n6905) );
  HS65_LS_NAND2X2 U12569 ( .A(n239), .B(n267), .Z(n5313) );
  HS65_LS_NAND2X2 U12570 ( .A(n458), .B(n486), .Z(n5428) );
  HS65_LS_NAND2X2 U12571 ( .A(n281), .B(n309), .Z(n7020) );
  HS65_LS_NAND2X2 U12572 ( .A(n683), .B(n705), .Z(n5197) );
  HS65_LS_NAND2X2 U12573 ( .A(n501), .B(n523), .Z(n6789) );
  HS65_LS_NAND2X2 U12574 ( .A(n457), .B(n486), .Z(n5405) );
  HS65_LS_NAND2X2 U12575 ( .A(n238), .B(n267), .Z(n5290) );
  HS65_LS_NAND2X2 U12576 ( .A(n684), .B(n705), .Z(n5173) );
  HS65_LS_NAND2X2 U12577 ( .A(n280), .B(n309), .Z(n6997) );
  HS65_LS_NAND2X2 U12578 ( .A(n59), .B(n88), .Z(n6882) );
  HS65_LS_NAND2X2 U12579 ( .A(n502), .B(n523), .Z(n6765) );
  HS65_LS_NOR4ABX2 U12580 ( .A(n6667), .B(n6668), .C(n6669), .D(n6670), .Z(
        n6660) );
  HS65_LS_NOR4ABX2 U12581 ( .A(n5074), .B(n5075), .C(n5076), .D(n5077), .Z(
        n5067) );
  HS65_LS_NAND2X2 U12582 ( .A(n358), .B(n336), .Z(n8358) );
  HS65_LS_NAND2X2 U12583 ( .A(n447), .B(n421), .Z(n3388) );
  HS65_LS_NAND2X2 U12584 ( .A(n430), .B(n411), .Z(n3195) );
  HS65_LS_NOR4ABX2 U12585 ( .A(n4210), .B(n3520), .C(n3109), .D(n3437), .Z(
        n4207) );
  HS65_LS_OAI21X2 U12586 ( .A(n194), .B(n192), .C(n212), .Z(n4210) );
  HS65_LS_NAND2X2 U12587 ( .A(n468), .B(n486), .Z(n4986) );
  HS65_LS_NAND2X2 U12588 ( .A(n249), .B(n267), .Z(n4932) );
  HS65_LS_NAND2X2 U12589 ( .A(n676), .B(n705), .Z(n4856) );
  HS65_LS_NAND2X2 U12590 ( .A(n291), .B(n309), .Z(n6579) );
  HS65_LS_NAND2X2 U12591 ( .A(n70), .B(n88), .Z(n6525) );
  HS65_LS_NAND2X2 U12592 ( .A(n494), .B(n523), .Z(n6449) );
  HS65_LS_NAND2X2 U12593 ( .A(n11), .B(n41), .Z(n4716) );
  HS65_LS_NAND2X2 U12594 ( .A(n537), .B(n567), .Z(n6309) );
  HS65_LS_NAND2X2 U12595 ( .A(n216), .B(n195), .Z(n3436) );
  HS65_LSS_XNOR2X3 U12596 ( .A(n3018), .B(n2771), .Z(n6004) );
  HS65_LSS_XNOR2X3 U12597 ( .A(n3222), .B(n2779), .Z(n4411) );
  HS65_LS_NAND4ABX3 U12598 ( .A(n2500), .B(n2266), .C(n2501), .D(n2502), .Z(
        n2499) );
  HS65_LS_NAND4ABX3 U12599 ( .A(n1748), .B(n1514), .C(n1749), .D(n1750), .Z(
        n1747) );
  HS65_LS_NAND2X2 U12600 ( .A(n121), .B(n107), .Z(n7921) );
  HS65_LS_NAND2X2 U12601 ( .A(n608), .B(n594), .Z(n7822) );
  HS65_LSS_XOR2X3 U12602 ( .A(n3217), .B(n2774), .Z(n5991) );
  HS65_LSS_XOR2X3 U12603 ( .A(n3225), .B(n2782), .Z(n4398) );
  HS65_LS_NOR4ABX2 U12604 ( .A(n8417), .B(n8761), .C(n8711), .D(n8427), .Z(
        n9026) );
  HS65_LS_NOR4ABX2 U12605 ( .A(n8477), .B(n8849), .C(n8799), .D(n8487), .Z(
        n9084) );
  HS65_LS_OAI21X2 U12606 ( .A(n200), .B(n3085), .C(n210), .Z(n3082) );
  HS65_LS_NAND2X2 U12607 ( .A(n417), .B(n439), .Z(n3878) );
  HS65_LS_OAI21X2 U12608 ( .A(n332), .B(n8346), .C(n341), .Z(n8343) );
  HS65_LS_NAND3AX3 U12609 ( .A(n2293), .B(n2294), .C(n2275), .Z(n2292) );
  HS65_LS_NAND3AX3 U12610 ( .A(n1541), .B(n1542), .C(n1523), .Z(n1540) );
  HS65_LS_NAND3AX3 U12611 ( .A(n1165), .B(n1166), .C(n1147), .Z(n1164) );
  HS65_LS_NAND3AX3 U12612 ( .A(n1917), .B(n1918), .C(n1899), .Z(n1916) );
  HS65_LS_NOR4ABX2 U12613 ( .A(n8253), .B(n8295), .C(n8219), .D(n8288), .Z(
        n8962) );
  HS65_LS_NAND2X2 U12614 ( .A(n378), .B(n387), .Z(n8211) );
  HS65_LS_NAND2X2 U12615 ( .A(n199), .B(n226), .Z(n3428) );
  HS65_LS_NOR4ABX2 U12616 ( .A(n3393), .B(n3848), .C(n3873), .D(n3866), .Z(
        n4329) );
  HS65_LS_NOR2X2 U12617 ( .A(n903), .B(n904), .Z(n2334) );
  HS65_LS_NOR2X2 U12618 ( .A(n821), .B(n822), .Z(n1582) );
  HS65_LS_NAND2X2 U12619 ( .A(n903), .B(n916), .Z(n2506) );
  HS65_LS_NAND2X2 U12620 ( .A(n821), .B(n834), .Z(n1754) );
  HS65_LS_NOR2X2 U12621 ( .A(n862), .B(n863), .Z(n1206) );
  HS65_LS_NOR2X2 U12622 ( .A(n780), .B(n781), .Z(n1958) );
  HS65_LS_OAI21X2 U12623 ( .A(n641), .B(n3314), .C(n662), .Z(n3311) );
  HS65_LS_NAND2X2 U12624 ( .A(n862), .B(n875), .Z(n1378) );
  HS65_LS_NOR4ABX2 U12625 ( .A(n3331), .B(n3756), .C(n3730), .D(n3749), .Z(
        n4270) );
  HS65_LS_OAI21X2 U12626 ( .A(n381), .B(n8093), .C(n403), .Z(n8102) );
  HS65_LS_NOR2X2 U12627 ( .A(n83), .B(n79), .Z(n6479) );
  HS65_LS_NOR2X2 U12628 ( .A(n304), .B(n300), .Z(n6593) );
  HS65_LS_NOR2X2 U12629 ( .A(n262), .B(n258), .Z(n4886) );
  HS65_LS_NOR2X2 U12630 ( .A(n481), .B(n477), .Z(n5000) );
  HS65_LS_NOR2X2 U12631 ( .A(n700), .B(n696), .Z(n4872) );
  HS65_LS_NOR2X2 U12632 ( .A(n518), .B(n514), .Z(n6465) );
  HS65_LS_NOR2X2 U12633 ( .A(n171), .B(n167), .Z(n3289) );
  HS65_LS_NOR2X2 U12634 ( .A(n439), .B(n435), .Z(n3413) );
  HS65_LS_NAND2X2 U12635 ( .A(n780), .B(n793), .Z(n2130) );
  HS65_LS_NOR2X2 U12636 ( .A(n36), .B(n32), .Z(n4668) );
  HS65_LS_NOR2X2 U12637 ( .A(n562), .B(n558), .Z(n6261) );
  HS65_LS_NAND2X2 U12638 ( .A(n612), .B(n583), .Z(n8761) );
  HS65_LS_NAND2X2 U12639 ( .A(n125), .B(n96), .Z(n8849) );
  HS65_LS_OAI21X2 U12640 ( .A(n372), .B(n365), .C(n404), .Z(n8664) );
  HS65_LS_NOR2X2 U12641 ( .A(n663), .B(n659), .Z(n3351) );
  HS65_LS_NOR2X2 U12642 ( .A(n218), .B(n213), .Z(n3125) );
  HS65_LS_NAND2X2 U12643 ( .A(n667), .B(n647), .Z(n3738) );
  HS65_LSS_XOR2X3 U12644 ( .A(n3221), .B(n2778), .Z(n4416) );
  HS65_LSS_XOR2X3 U12645 ( .A(n3017), .B(n2770), .Z(n6009) );
  HS65_LS_NAND2X2 U12646 ( .A(n218), .B(n198), .Z(n3539) );
  HS65_LS_NAND2X2 U12647 ( .A(n901), .B(n919), .Z(n2450) );
  HS65_LS_NAND2X2 U12648 ( .A(n819), .B(n837), .Z(n1698) );
  HS65_LS_NAND2X2 U12649 ( .A(n860), .B(n878), .Z(n1322) );
  HS65_LS_NAND2X2 U12650 ( .A(n778), .B(n796), .Z(n2074) );
  HS65_LS_NAND2X2 U12651 ( .A(n219), .B(n192), .Z(n3496) );
  HS65_LS_NAND2X2 U12652 ( .A(n227), .B(n205), .Z(n2952) );
  HS65_LS_NAND2X2 U12653 ( .A(n439), .B(n414), .Z(n3896) );
  HS65_LS_NAND2X2 U12654 ( .A(n443), .B(n423), .Z(n3855) );
  HS65_LSS_XOR2X3 U12655 ( .A(n2810), .B(n2786), .Z(n2628) );
  HS65_LS_NAND2X2 U12656 ( .A(n654), .B(n634), .Z(n3154) );
  HS65_LS_OAI21X2 U12657 ( .A(n417), .B(n3376), .C(n438), .Z(n3373) );
  HS65_LSS_XOR2X3 U12658 ( .A(n2826), .B(n2802), .Z(n4382) );
  HS65_LS_NOR2X2 U12659 ( .A(n420), .B(n3787), .Z(n3842) );
  HS65_LS_NAND4ABX3 U12660 ( .A(n2348), .B(n2349), .C(n2350), .D(n2351), .Z(
        n2293) );
  HS65_LS_NAND4ABX3 U12661 ( .A(n2377), .B(n2378), .C(n2379), .D(n2380), .Z(
        n2349) );
  HS65_LS_NOR4ABX2 U12662 ( .A(n2352), .B(n2353), .C(n2354), .D(n2355), .Z(
        n2351) );
  HS65_LS_MX41X4 U12663 ( .D0(n919), .S0(n900), .D1(n930), .S1(n897), .D2(n915), .S2(n905), .D3(n927), .S3(n901), .Z(n2348) );
  HS65_LS_NAND4ABX3 U12664 ( .A(n1596), .B(n1597), .C(n1598), .D(n1599), .Z(
        n1541) );
  HS65_LS_NAND4ABX3 U12665 ( .A(n1625), .B(n1626), .C(n1627), .D(n1628), .Z(
        n1597) );
  HS65_LS_NOR4ABX2 U12666 ( .A(n1600), .B(n1601), .C(n1602), .D(n1603), .Z(
        n1599) );
  HS65_LS_MX41X4 U12667 ( .D0(n837), .S0(n818), .D1(n848), .S1(n815), .D2(n833), .S2(n823), .D3(n845), .S3(n819), .Z(n1596) );
  HS65_LS_NAND4ABX3 U12668 ( .A(n1220), .B(n1221), .C(n1222), .D(n1223), .Z(
        n1165) );
  HS65_LS_NAND4ABX3 U12669 ( .A(n1249), .B(n1250), .C(n1251), .D(n1252), .Z(
        n1221) );
  HS65_LS_NOR4ABX2 U12670 ( .A(n1224), .B(n1225), .C(n1226), .D(n1227), .Z(
        n1223) );
  HS65_LS_MX41X4 U12671 ( .D0(n878), .S0(n859), .D1(n889), .S1(n856), .D2(n874), .S2(n864), .D3(n886), .S3(n860), .Z(n1220) );
  HS65_LS_NAND4ABX3 U12672 ( .A(n1972), .B(n1973), .C(n1974), .D(n1975), .Z(
        n1917) );
  HS65_LS_NAND4ABX3 U12673 ( .A(n2001), .B(n2002), .C(n2003), .D(n2004), .Z(
        n1973) );
  HS65_LS_NOR4ABX2 U12674 ( .A(n1976), .B(n1977), .C(n1978), .D(n1979), .Z(
        n1975) );
  HS65_LS_MX41X4 U12675 ( .D0(n796), .S0(n777), .D1(n807), .S1(n774), .D2(n792), .S2(n782), .D3(n804), .S3(n778), .Z(n1972) );
  HS65_LS_OAI21X2 U12676 ( .A(n155), .B(n3247), .C(n165), .Z(n3244) );
  HS65_LS_OAI21X2 U12677 ( .A(n921), .B(n2356), .C(n895), .Z(n2353) );
  HS65_LS_OAI21X2 U12678 ( .A(n839), .B(n1604), .C(n813), .Z(n1601) );
  HS65_LS_NOR2X2 U12679 ( .A(n542), .B(n6607), .Z(n6631) );
  HS65_LS_NOR2X2 U12680 ( .A(n16), .B(n5014), .Z(n5038) );
  HS65_LS_NOR2X2 U12681 ( .A(n64), .B(n6846), .Z(n6869) );
  HS65_LS_NOR2X2 U12682 ( .A(n243), .B(n5254), .Z(n5277) );
  HS65_LS_NOR2X2 U12683 ( .A(n462), .B(n5369), .Z(n5392) );
  HS65_LS_NOR2X2 U12684 ( .A(n285), .B(n6961), .Z(n6984) );
  HS65_LS_NOR2X2 U12685 ( .A(n681), .B(n5136), .Z(n5160) );
  HS65_LS_NOR2X2 U12686 ( .A(n499), .B(n6728), .Z(n6752) );
  HS65_LS_OAI21X2 U12687 ( .A(n880), .B(n1228), .C(n854), .Z(n1225) );
  HS65_LS_OAI21X2 U12688 ( .A(n798), .B(n1980), .C(n772), .Z(n1977) );
  HS65_LS_NAND2X2 U12689 ( .A(n326), .B(n346), .Z(n8562) );
  HS65_LS_NAND2X2 U12690 ( .A(n919), .B(n896), .Z(n2311) );
  HS65_LS_NAND2X2 U12691 ( .A(n837), .B(n814), .Z(n1559) );
  HS65_LS_IVX2 U12692 ( .A(n2701), .Z(n409) );
  HS65_LS_NAND2X2 U12693 ( .A(n622), .B(n598), .Z(n8724) );
  HS65_LS_NAND2X2 U12694 ( .A(n135), .B(n111), .Z(n8812) );
  HS65_LS_NAND2X2 U12695 ( .A(n878), .B(n855), .Z(n1183) );
  HS65_LS_NAND2X2 U12696 ( .A(n796), .B(n773), .Z(n1935) );
  HS65_LS_NAND4ABX3 U12697 ( .A(n3923), .B(n3924), .C(n3925), .D(n3926), .Z(
        n3917) );
  HS65_LS_AOI212X2 U12698 ( .A(n148), .B(n180), .C(n181), .D(n144), .E(n3927), 
        .Z(n3926) );
  HS65_LS_NAND2X2 U12699 ( .A(n167), .B(n152), .Z(n3638) );
  HS65_LS_NAND2X2 U12700 ( .A(n423), .B(n442), .Z(n3199) );
  HS65_LS_NAND2X2 U12701 ( .A(n192), .B(n215), .Z(n2956) );
  HS65_LS_NAND2X2 U12702 ( .A(n647), .B(n666), .Z(n3158) );
  HS65_LS_NAND2X2 U12703 ( .A(n394), .B(n380), .Z(n8298) );
  HS65_LS_NAND2X2 U12704 ( .A(n356), .B(n331), .Z(n8602) );
  HS65_LS_NAND4ABX3 U12705 ( .A(n4538), .B(n4539), .C(n4540), .D(n4541), .Z(
        n4528) );
  HS65_LS_AOI212X2 U12706 ( .A(n680), .B(n697), .C(n676), .D(n712), .E(n4542), 
        .Z(n4541) );
  HS65_LS_NAND4ABX3 U12707 ( .A(n6189), .B(n6190), .C(n6191), .D(n6192), .Z(
        n6181) );
  HS65_LS_AOI212X2 U12708 ( .A(n66), .B(n80), .C(n70), .D(n74), .E(n6193), .Z(
        n6192) );
  HS65_LS_NAND4ABX3 U12709 ( .A(n6131), .B(n6132), .C(n6133), .D(n6134), .Z(
        n6121) );
  HS65_LS_AOI212X2 U12710 ( .A(n498), .B(n515), .C(n494), .D(n530), .E(n6135), 
        .Z(n6134) );
  HS65_LS_NAND4ABX3 U12711 ( .A(n4596), .B(n4597), .C(n4598), .D(n4599), .Z(
        n4588) );
  HS65_LS_AOI212X2 U12712 ( .A(n245), .B(n259), .C(n249), .D(n253), .E(n4600), 
        .Z(n4599) );
  HS65_LS_NAND2X2 U12713 ( .A(n647), .B(n660), .Z(n3326) );
  HS65_LSS_XOR3X2 U12714 ( .A(n2674), .B(n2637), .C(n2711), .Z(n2749) );
  HS65_LSS_XNOR3X2 U12715 ( .A(n2667), .B(n2661), .C(n2666), .Z(n2665) );
  HS65_LS_NAND2X2 U12716 ( .A(n663), .B(n637), .Z(n3779) );
  HS65_LS_NAND2X2 U12717 ( .A(n478), .B(n453), .Z(n5386) );
  HS65_LS_NAND2X2 U12718 ( .A(n259), .B(n234), .Z(n5271) );
  HS65_LS_NAND2X2 U12719 ( .A(n697), .B(n687), .Z(n5154) );
  HS65_LS_NAND2X2 U12720 ( .A(n301), .B(n276), .Z(n6978) );
  HS65_LS_NAND2X2 U12721 ( .A(n80), .B(n55), .Z(n6863) );
  HS65_LS_NAND2X2 U12722 ( .A(n515), .B(n505), .Z(n6746) );
  HS65_LS_OAI21X2 U12723 ( .A(n422), .B(n423), .C(n437), .Z(n4327) );
  HS65_LS_NAND2X2 U12724 ( .A(n331), .B(n352), .Z(n8544) );
  HS65_LS_NAND2X2 U12725 ( .A(n599), .B(n619), .Z(n7806) );
  HS65_LS_NAND2X2 U12726 ( .A(n112), .B(n132), .Z(n7906) );
  HS65_LS_OAI21X2 U12727 ( .A(n795), .B(n796), .C(n786), .Z(n2229) );
  HS65_LS_OAI21X2 U12728 ( .A(n877), .B(n878), .C(n868), .Z(n1477) );
  HS65_LS_NAND2X2 U12729 ( .A(n670), .B(n637), .Z(n3761) );
  HS65_LS_IVX2 U12730 ( .A(n2717), .Z(n408) );
  HS65_LS_NAND2X2 U12731 ( .A(n143), .B(n168), .Z(n3639) );
  HS65_LS_NAND2X2 U12732 ( .A(n77), .B(n66), .Z(n6866) );
  HS65_LS_NAND2X2 U12733 ( .A(n256), .B(n245), .Z(n5274) );
  HS65_LS_NAND2X2 U12734 ( .A(n475), .B(n464), .Z(n5389) );
  HS65_LS_NAND2X2 U12735 ( .A(n298), .B(n287), .Z(n6981) );
  HS65_LS_NAND2X2 U12736 ( .A(n709), .B(n680), .Z(n5157) );
  HS65_LS_NAND2X2 U12737 ( .A(n527), .B(n498), .Z(n6749) );
  HS65_LS_NAND2X2 U12738 ( .A(n42), .B(n25), .Z(n5111) );
  HS65_LS_NAND2X2 U12739 ( .A(n568), .B(n551), .Z(n6704) );
  HS65_LS_AOI12X2 U12740 ( .A(n613), .B(n583), .C(n8758), .Z(n8755) );
  HS65_LS_AOI12X2 U12741 ( .A(n126), .B(n96), .C(n8846), .Z(n8843) );
  HS65_LS_NOR2X2 U12742 ( .A(n615), .B(n625), .Z(n8430) );
  HS65_LS_NOR2X2 U12743 ( .A(n128), .B(n138), .Z(n8441) );
  HS65_LS_IVX2 U12744 ( .A(n2669), .Z(n141) );
  HS65_LS_NAND2X2 U12745 ( .A(n335), .B(n350), .Z(n8381) );
  HS65_LS_NAND3AX3 U12746 ( .A(n8210), .B(n8211), .C(n8212), .Z(n8209) );
  HS65_LS_NAND2X2 U12747 ( .A(n324), .B(n346), .Z(n8603) );
  HS65_LS_NAND2X2 U12748 ( .A(n606), .B(n584), .Z(n8695) );
  HS65_LS_NAND2X2 U12749 ( .A(n119), .B(n97), .Z(n8783) );
  HS65_LS_NAND3AX3 U12750 ( .A(n6848), .B(n6849), .C(n6850), .Z(n6847) );
  HS65_LS_NAND3AX3 U12751 ( .A(n5256), .B(n5257), .C(n5258), .Z(n5255) );
  HS65_LS_NAND3AX3 U12752 ( .A(n5371), .B(n5372), .C(n5373), .Z(n5370) );
  HS65_LS_NAND3AX3 U12753 ( .A(n6963), .B(n6964), .C(n6965), .Z(n6962) );
  HS65_LS_NAND3AX3 U12754 ( .A(n6730), .B(n6731), .C(n6732), .Z(n6729) );
  HS65_LS_NAND3AX3 U12755 ( .A(n5138), .B(n5139), .C(n5140), .Z(n5137) );
  HS65_LS_NAND2X2 U12756 ( .A(n156), .B(n170), .Z(n3039) );
  HS65_LS_NAND2X2 U12757 ( .A(n321), .B(n357), .Z(n8566) );
  HS65_LSS_XOR3X2 U12758 ( .A(n7556), .B(n2628), .C(n2762), .Z(n7569) );
  HS65_LS_NAND2X2 U12759 ( .A(n366), .B(n393), .Z(n8262) );
  HS65_LS_NOR2X2 U12760 ( .A(n399), .B(n402), .Z(n8129) );
  HS65_LS_NAND2X2 U12761 ( .A(n147), .B(n176), .Z(n3283) );
  HS65_LS_NAND2X2 U12762 ( .A(n147), .B(n175), .Z(n3254) );
  HS65_LS_NAND3AX3 U12763 ( .A(n6609), .B(n6610), .C(n6611), .Z(n6608) );
  HS65_LS_NAND3AX3 U12764 ( .A(n5016), .B(n5017), .C(n5018), .Z(n5015) );
  HS65_LS_NAND2X2 U12765 ( .A(n840), .B(n826), .Z(n1678) );
  HS65_LS_NAND2X2 U12766 ( .A(n922), .B(n908), .Z(n2430) );
  HS65_LS_NAND2X2 U12767 ( .A(n881), .B(n867), .Z(n1302) );
  HS65_LS_NOR2X2 U12768 ( .A(n925), .B(n922), .Z(n2503) );
  HS65_LS_NOR2X2 U12769 ( .A(n843), .B(n840), .Z(n1751) );
  HS65_LS_NAND2X2 U12770 ( .A(n799), .B(n785), .Z(n2054) );
  HS65_LS_NOR2X2 U12771 ( .A(n884), .B(n881), .Z(n1375) );
  HS65_LS_NOR2X2 U12772 ( .A(n802), .B(n799), .Z(n2127) );
  HS65_LS_NOR2X2 U12773 ( .A(n927), .B(n916), .Z(n2391) );
  HS65_LS_NOR2X2 U12774 ( .A(n845), .B(n834), .Z(n1639) );
  HS65_LS_NOR2X2 U12775 ( .A(n886), .B(n875), .Z(n1263) );
  HS65_LS_NOR2X2 U12776 ( .A(n804), .B(n793), .Z(n2015) );
  HS65_LS_NOR2X2 U12777 ( .A(n201), .B(n204), .Z(n3535) );
  HS65_LS_NOR2X2 U12778 ( .A(n640), .B(n636), .Z(n3775) );
  HS65_LS_NOR2X2 U12779 ( .A(n329), .B(n331), .Z(n8378) );
  HS65_LS_NOR2X2 U12780 ( .A(n416), .B(n413), .Z(n3892) );
  HS65_LS_NOR2X2 U12781 ( .A(n379), .B(n377), .Z(n8314) );
  HS65_LS_NAND2X2 U12782 ( .A(n413), .B(n431), .Z(n3835) );
  HS65_LS_NOR2X2 U12783 ( .A(n639), .B(n637), .Z(n3349) );
  HS65_LS_NAND2X2 U12784 ( .A(n612), .B(n598), .Z(n8709) );
  HS65_LS_NAND2X2 U12785 ( .A(n125), .B(n111), .Z(n8797) );
  HS65_LS_NAND2X2 U12786 ( .A(n204), .B(n228), .Z(n3476) );
  HS65_LS_NAND2X2 U12787 ( .A(n636), .B(n655), .Z(n3719) );
  HS65_LS_NAND2X2 U12788 ( .A(n354), .B(n326), .Z(n8601) );
  HS65_LS_NAND2X2 U12789 ( .A(n106), .B(n124), .Z(n7937) );
  HS65_LS_NAND2X2 U12790 ( .A(n593), .B(n611), .Z(n7838) );
  HS65_LS_NAND2X2 U12791 ( .A(n482), .B(n460), .Z(n5477) );
  HS65_LS_NAND2X2 U12792 ( .A(n263), .B(n241), .Z(n5362) );
  HS65_LS_NAND2X2 U12793 ( .A(n702), .B(n686), .Z(n5247) );
  HS65_LS_NAND2X2 U12794 ( .A(n305), .B(n283), .Z(n7069) );
  HS65_LS_NAND2X2 U12795 ( .A(n84), .B(n62), .Z(n6954) );
  HS65_LS_NAND2X2 U12796 ( .A(n520), .B(n504), .Z(n6839) );
  HS65_LS_NOR2X2 U12797 ( .A(n154), .B(n153), .Z(n3278) );
  HS65_LS_NAND2X2 U12798 ( .A(n865), .B(n880), .Z(n1279) );
  HS65_LS_NAND2X2 U12799 ( .A(n783), .B(n798), .Z(n2031) );
  HS65_LS_NAND2X2 U12800 ( .A(n906), .B(n921), .Z(n2407) );
  HS65_LS_NAND2X2 U12801 ( .A(n824), .B(n839), .Z(n1655) );
  HS65_LS_OAI21X2 U12802 ( .A(n586), .B(n8400), .C(n611), .Z(n8425) );
  HS65_LS_OAI21X2 U12803 ( .A(n99), .B(n8460), .C(n124), .Z(n8485) );
  HS65_LS_NAND2X2 U12804 ( .A(n904), .B(n916), .Z(n2477) );
  HS65_LS_NAND2X2 U12805 ( .A(n822), .B(n834), .Z(n1725) );
  HS65_LS_OAI21X2 U12806 ( .A(n334), .B(n318), .C(n345), .Z(n8872) );
  HS65_LS_NAND2X2 U12807 ( .A(n863), .B(n875), .Z(n1349) );
  HS65_LS_NAND2X2 U12808 ( .A(n781), .B(n793), .Z(n2101) );
  HS65_LS_MX41X4 U12809 ( .D0(n584), .S0(n618), .D1(n608), .S1(n600), .D2(n623), .S2(n586), .D3(n612), .S3(n599), .Z(n8756) );
  HS65_LS_MX41X4 U12810 ( .D0(n97), .S0(n131), .D1(n121), .S1(n113), .D2(n136), 
        .S2(n99), .D3(n125), .S3(n112), .Z(n8844) );
  HS65_LS_NAND2X2 U12811 ( .A(n435), .B(n414), .Z(n3882) );
  HS65_LS_NAND4ABX3 U12812 ( .A(n1661), .B(n1756), .C(n1829), .D(n1637), .Z(
        n1825) );
  HS65_LS_OAI21X2 U12813 ( .A(n846), .B(n838), .C(n823), .Z(n1829) );
  HS65_LS_NAND4ABX3 U12814 ( .A(n2413), .B(n2508), .C(n2581), .D(n2389), .Z(
        n2577) );
  HS65_LS_OAI21X2 U12815 ( .A(n928), .B(n920), .C(n905), .Z(n2581) );
  HS65_LS_NAND4ABX3 U12816 ( .A(n1285), .B(n1380), .C(n1453), .D(n1261), .Z(
        n1449) );
  HS65_LS_OAI21X2 U12817 ( .A(n887), .B(n879), .C(n864), .Z(n1453) );
  HS65_LS_NAND4ABX3 U12818 ( .A(n2037), .B(n2132), .C(n2205), .D(n2013), .Z(
        n2201) );
  HS65_LS_OAI21X2 U12819 ( .A(n805), .B(n797), .C(n782), .Z(n2205) );
  HS65_LS_NAND4ABX3 U12820 ( .A(n3802), .B(n3898), .C(n4316), .D(n3409), .Z(
        n4312) );
  HS65_LS_OAI21X2 U12821 ( .A(n421), .B(n419), .C(n434), .Z(n4316) );
  HS65_LS_NAND4ABX3 U12822 ( .A(n3685), .B(n3781), .C(n4257), .D(n3347), .Z(
        n4253) );
  HS65_LS_OAI21X2 U12823 ( .A(n645), .B(n643), .C(n658), .Z(n4257) );
  HS65_LS_NAND4ABX3 U12824 ( .A(n6635), .B(n6636), .C(n6637), .D(n6638), .Z(
        n6620) );
  HS65_LS_NAND4ABX3 U12825 ( .A(n5042), .B(n5043), .C(n5044), .D(n5045), .Z(
        n5027) );
  HS65_LS_NAND2X2 U12826 ( .A(n919), .B(n898), .Z(n2308) );
  HS65_LS_NAND2X2 U12827 ( .A(n837), .B(n816), .Z(n1556) );
  HS65_LS_NAND4ABX3 U12828 ( .A(n6873), .B(n6874), .C(n6875), .D(n6876), .Z(
        n6858) );
  HS65_LS_NAND4ABX3 U12829 ( .A(n5281), .B(n5282), .C(n5283), .D(n5284), .Z(
        n5266) );
  HS65_LS_NAND4ABX3 U12830 ( .A(n5396), .B(n5397), .C(n5398), .D(n5399), .Z(
        n5381) );
  HS65_LS_NAND4ABX3 U12831 ( .A(n6988), .B(n6989), .C(n6990), .D(n6991), .Z(
        n6973) );
  HS65_LS_NAND4ABX3 U12832 ( .A(n5164), .B(n5165), .C(n5166), .D(n5167), .Z(
        n5149) );
  HS65_LS_NAND4ABX3 U12833 ( .A(n6756), .B(n6757), .C(n6758), .D(n6759), .Z(
        n6741) );
  HS65_LS_NAND2X2 U12834 ( .A(n878), .B(n857), .Z(n1180) );
  HS65_LS_NAND2X2 U12835 ( .A(n796), .B(n775), .Z(n1932) );
  HS65_LS_NAND4ABX3 U12836 ( .A(n8221), .B(n8222), .C(n8223), .D(n8224), .Z(
        n8214) );
  HS65_LS_NAND4ABX3 U12837 ( .A(n3507), .B(n3508), .C(n3509), .D(n3510), .Z(
        n3491) );
  HS65_LS_NAND4ABX3 U12838 ( .A(n3748), .B(n3749), .C(n3750), .D(n3751), .Z(
        n3733) );
  HS65_LS_NAND4ABX3 U12839 ( .A(n2456), .B(n2457), .C(n2458), .D(n2459), .Z(
        n2446) );
  HS65_LS_NAND4ABX3 U12840 ( .A(n1704), .B(n1705), .C(n1706), .D(n1707), .Z(
        n1694) );
  HS65_LS_NAND4ABX3 U12841 ( .A(n1328), .B(n1329), .C(n1330), .D(n1331), .Z(
        n1318) );
  HS65_LS_NAND4ABX3 U12842 ( .A(n2080), .B(n2081), .C(n2082), .D(n2083), .Z(
        n2070) );
  HS65_LS_NAND3AX3 U12843 ( .A(n3346), .B(n3347), .C(n3348), .Z(n3340) );
  HS65_LS_OAI21X2 U12844 ( .A(n645), .B(n3314), .C(n654), .Z(n3348) );
  HS65_LS_NAND2X2 U12845 ( .A(n370), .B(n397), .Z(n8087) );
  HS65_LS_NAND3AX3 U12846 ( .A(n2388), .B(n2389), .C(n2390), .Z(n2382) );
  HS65_LS_OAI21X2 U12847 ( .A(n928), .B(n2356), .C(n898), .Z(n2390) );
  HS65_LS_NAND3AX3 U12848 ( .A(n1636), .B(n1637), .C(n1638), .Z(n1630) );
  HS65_LS_OAI21X2 U12849 ( .A(n846), .B(n1604), .C(n816), .Z(n1638) );
  HS65_LS_NAND3AX3 U12850 ( .A(n1260), .B(n1261), .C(n1262), .Z(n1254) );
  HS65_LS_OAI21X2 U12851 ( .A(n887), .B(n1228), .C(n857), .Z(n1262) );
  HS65_LS_NAND3AX3 U12852 ( .A(n2012), .B(n2013), .C(n2014), .Z(n2006) );
  HS65_LS_OAI21X2 U12853 ( .A(n805), .B(n1980), .C(n775), .Z(n2014) );
  HS65_LS_NAND4ABX3 U12854 ( .A(n3846), .B(n3847), .C(n3848), .D(n3849), .Z(
        n3831) );
  HS65_LS_NAND3AX3 U12855 ( .A(n3103), .B(n3104), .C(n3105), .Z(n3088) );
  HS65_LS_AOI12X2 U12856 ( .A(n189), .B(n3106), .C(n3107), .Z(n3105) );
  HS65_LS_NAND3AX3 U12857 ( .A(n3265), .B(n3266), .C(n3267), .Z(n3250) );
  HS65_LS_AOI12X2 U12858 ( .A(n143), .B(n3268), .C(n3269), .Z(n3267) );
  HS65_LS_NAND3AX3 U12859 ( .A(n1244), .B(n1245), .C(n1246), .Z(n1231) );
  HS65_LS_AOI12X2 U12860 ( .A(n882), .B(n1247), .C(n1248), .Z(n1246) );
  HS65_LS_NAND3AX3 U12861 ( .A(n1996), .B(n1997), .C(n1998), .Z(n1983) );
  HS65_LS_AOI12X2 U12862 ( .A(n800), .B(n1999), .C(n2000), .Z(n1998) );
  HS65_LS_NAND3AX3 U12863 ( .A(n3392), .B(n3393), .C(n3394), .Z(n3379) );
  HS65_LS_AOI12X2 U12864 ( .A(n424), .B(n3395), .C(n3396), .Z(n3394) );
  HS65_LS_NAND4ABX3 U12865 ( .A(n8424), .B(n8416), .C(n8749), .D(n9036), .Z(
        n9032) );
  HS65_LS_OAI21X2 U12866 ( .A(n618), .B(n614), .C(n592), .Z(n9036) );
  HS65_LS_NAND4ABX3 U12867 ( .A(n8484), .B(n8476), .C(n8837), .D(n9094), .Z(
        n9090) );
  HS65_LS_OAI21X2 U12868 ( .A(n131), .B(n127), .C(n105), .Z(n9094) );
  HS65_LS_NAND3AX3 U12869 ( .A(n7824), .B(n8413), .C(n8414), .Z(n8403) );
  HS65_LS_AOI12X2 U12870 ( .A(n591), .B(n7841), .C(n8415), .Z(n8414) );
  HS65_LS_NAND3AX3 U12871 ( .A(n7923), .B(n8473), .C(n8474), .Z(n8463) );
  HS65_LS_AOI12X2 U12872 ( .A(n104), .B(n7940), .C(n8475), .Z(n8474) );
  HS65_LS_AOI12X2 U12873 ( .A(n398), .B(n371), .C(n8232), .Z(n8229) );
  HS65_LS_NAND4ABX3 U12874 ( .A(n3406), .B(n3823), .C(n3890), .D(n3383), .Z(
        n4324) );
  HS65_LS_NAND4ABX3 U12875 ( .A(n3861), .B(n3862), .C(n3863), .D(n3864), .Z(
        n3851) );
  HS65_LS_AOI12X2 U12876 ( .A(n169), .B(n153), .C(n3555), .Z(n4159) );
  HS65_LS_NAND3X2 U12877 ( .A(n6530), .B(n6531), .C(n6532), .Z(n6516) );
  HS65_LS_AOI12X2 U12878 ( .A(n68), .B(n6533), .C(n6534), .Z(n6532) );
  HS65_LS_NAND3X2 U12879 ( .A(n6584), .B(n6585), .C(n6586), .Z(n6570) );
  HS65_LS_AOI12X2 U12880 ( .A(n289), .B(n6587), .C(n6588), .Z(n6586) );
  HS65_LS_NAND3X2 U12881 ( .A(n4991), .B(n4992), .C(n4993), .Z(n4977) );
  HS65_LS_AOI12X2 U12882 ( .A(n466), .B(n4994), .C(n4995), .Z(n4993) );
  HS65_LS_NAND3X2 U12883 ( .A(n4937), .B(n4938), .C(n4939), .Z(n4923) );
  HS65_LS_AOI12X2 U12884 ( .A(n247), .B(n4940), .C(n4941), .Z(n4939) );
  HS65_LS_NAND3X2 U12885 ( .A(n4863), .B(n4864), .C(n4865), .Z(n4847) );
  HS65_LS_AOI12X2 U12886 ( .A(n675), .B(n4866), .C(n4867), .Z(n4865) );
  HS65_LS_NAND3X2 U12887 ( .A(n6456), .B(n6457), .C(n6458), .Z(n6440) );
  HS65_LS_AOI12X2 U12888 ( .A(n493), .B(n6459), .C(n6460), .Z(n6458) );
  HS65_LS_IVX2 U12889 ( .A(n8078), .Z(n392) );
  HS65_LS_AOI12X2 U12890 ( .A(n921), .B(n905), .C(n2455), .Z(n2452) );
  HS65_LS_AOI12X2 U12891 ( .A(n839), .B(n823), .C(n1703), .Z(n1700) );
  HS65_LS_AOI12X2 U12892 ( .A(n880), .B(n864), .C(n1327), .Z(n1324) );
  HS65_LS_AOI12X2 U12893 ( .A(n798), .B(n782), .C(n2079), .Z(n2076) );
  HS65_LS_IVX2 U12894 ( .A(n3234), .Z(n173) );
  HS65_LS_IVX2 U12895 ( .A(n8388), .Z(n617) );
  HS65_LS_IVX2 U12896 ( .A(n8448), .Z(n130) );
  HS65_LS_AOI12X2 U12897 ( .A(n417), .B(n434), .C(n3860), .Z(n3857) );
  HS65_LS_IVX2 U12898 ( .A(n4678), .Z(n39) );
  HS65_LS_IVX2 U12899 ( .A(n6271), .Z(n565) );
  HS65_LS_AO212X4 U12900 ( .A(n924), .B(n2484), .C(n925), .D(n906), .E(n2611), 
        .Z(n2610) );
  HS65_LS_CB4I6X4 U12901 ( .A(n926), .B(n927), .C(n905), .D(n2509), .Z(n2611)
         );
  HS65_LS_AO212X4 U12902 ( .A(n842), .B(n1732), .C(n843), .D(n824), .E(n1859), 
        .Z(n1858) );
  HS65_LS_CB4I6X4 U12903 ( .A(n844), .B(n845), .C(n823), .D(n1757), .Z(n1859)
         );
  HS65_LS_AO212X4 U12904 ( .A(n883), .B(n1356), .C(n884), .D(n865), .E(n1483), 
        .Z(n1482) );
  HS65_LS_CB4I6X4 U12905 ( .A(n885), .B(n886), .C(n864), .D(n1381), .Z(n1483)
         );
  HS65_LS_AO212X4 U12906 ( .A(n801), .B(n2108), .C(n802), .D(n783), .E(n2235), 
        .Z(n2234) );
  HS65_LS_CB4I6X4 U12907 ( .A(n803), .B(n804), .C(n782), .D(n2133), .Z(n2235)
         );
  HS65_LS_AOI12X2 U12908 ( .A(n641), .B(n658), .C(n3743), .Z(n3740) );
  HS65_LS_AOI12X2 U12909 ( .A(n200), .B(n225), .C(n3502), .Z(n3499) );
  HS65_LS_IVX2 U12910 ( .A(n4950), .Z(n488) );
  HS65_LS_IVX2 U12911 ( .A(n4896), .Z(n269) );
  HS65_LS_IVX2 U12912 ( .A(n6543), .Z(n311) );
  HS65_LS_IVX2 U12913 ( .A(n4818), .Z(n703) );
  HS65_LS_IVX2 U12914 ( .A(n6411), .Z(n521) );
  HS65_LS_IVX2 U12915 ( .A(n6489), .Z(n90) );
  HS65_LS_NAND4ABX3 U12916 ( .A(n8683), .B(n8165), .C(n8434), .D(n8710), .Z(
        n9018) );
  HS65_LS_NAND4ABX3 U12917 ( .A(n8771), .B(n8197), .C(n8445), .D(n8798), .Z(
        n9076) );
  HS65_LS_NAND4ABX3 U12918 ( .A(n6484), .B(n6360), .C(n6849), .D(n6886), .Z(
        n7461) );
  HS65_LS_NAND4ABX3 U12919 ( .A(n5005), .B(n4806), .C(n5372), .D(n5409), .Z(
        n5928) );
  HS65_LS_NAND4ABX3 U12920 ( .A(n6598), .B(n6399), .C(n6964), .D(n7001), .Z(
        n7520) );
  HS65_LS_NAND4ABX3 U12921 ( .A(n4891), .B(n4767), .C(n5257), .D(n5294), .Z(
        n5869) );
  HS65_LS_NAND4ABX3 U12922 ( .A(n4877), .B(n4660), .C(n5139), .D(n5177), .Z(
        n5797) );
  HS65_LS_NAND4ABX3 U12923 ( .A(n6470), .B(n6253), .C(n6731), .D(n6769), .Z(
        n7389) );
  HS65_LS_NAND4ABX3 U12924 ( .A(n6266), .B(n6176), .C(n6610), .D(n6648), .Z(
        n7327) );
  HS65_LS_NAND4ABX3 U12925 ( .A(n4673), .B(n4583), .C(n5017), .D(n5055), .Z(
        n5735) );
  HS65_LS_IVX2 U12926 ( .A(n3072), .Z(n220) );
  HS65_LS_IVX2 U12927 ( .A(n3364), .Z(n444) );
  HS65_LS_IVX2 U12928 ( .A(n3710), .Z(n657) );
  HS65_LS_IVX2 U12929 ( .A(n3302), .Z(n668) );
  HS65_LS_AND4X3 U12930 ( .A(n1853), .B(n1628), .C(n1721), .D(n1655), .Z(n1847) );
  HS65_LS_OAI21X2 U12931 ( .A(n836), .B(n837), .C(n827), .Z(n1853) );
  HS65_LS_AND4X3 U12932 ( .A(n2605), .B(n2380), .C(n2473), .D(n2407), .Z(n2599) );
  HS65_LS_OAI21X2 U12933 ( .A(n918), .B(n919), .C(n909), .Z(n2605) );
  HS65_LS_IVX2 U12934 ( .A(n1593), .Z(n820) );
  HS65_LS_IVX2 U12935 ( .A(n2345), .Z(n902) );
  HS65_LS_IVX2 U12936 ( .A(n1969), .Z(n779) );
  HS65_LS_IVX2 U12937 ( .A(n1217), .Z(n861) );
  HS65_LS_NAND2X2 U12938 ( .A(n329), .B(n347), .Z(n8515) );
  HS65_LS_IVX2 U12939 ( .A(n8333), .Z(n355) );
  HS65_LS_IVX2 U12940 ( .A(n7815), .Z(n607) );
  HS65_LS_IVX2 U12941 ( .A(n7915), .Z(n120) );
  HS65_LS_IVX2 U12942 ( .A(n5439), .Z(n476) );
  HS65_LS_IVX2 U12943 ( .A(n7031), .Z(n299) );
  HS65_LS_IVX2 U12944 ( .A(n6916), .Z(n78) );
  HS65_LS_IVX2 U12945 ( .A(n5324), .Z(n257) );
  HS65_LS_IVX2 U12946 ( .A(n3827), .Z(n433) );
  HS65_LS_MX41X4 U12947 ( .D0(n919), .S0(n903), .D1(n923), .S1(n904), .D2(n920), .S2(n898), .D3(n915), .S3(n899), .Z(n2560) );
  HS65_LS_MX41X4 U12948 ( .D0(n837), .S0(n821), .D1(n841), .S1(n822), .D2(n838), .S2(n816), .D3(n833), .S3(n817), .Z(n1808) );
  HS65_LS_MX41X4 U12949 ( .D0(n796), .S0(n780), .D1(n800), .S1(n781), .D2(n797), .S2(n775), .D3(n792), .S3(n776), .Z(n2184) );
  HS65_LS_MX41X4 U12950 ( .D0(n878), .S0(n862), .D1(n882), .S1(n863), .D2(n879), .S2(n857), .D3(n874), .S3(n858), .Z(n1432) );
  HS65_LS_MX41X4 U12951 ( .D0(n366), .S0(n403), .D1(n395), .S1(n379), .D2(n380), .S2(n391), .D3(n378), .S3(n397), .Z(n8500) );
  HS65_LS_MX41X4 U12952 ( .D0(n920), .S0(n898), .D1(n922), .S1(n905), .D2(n915), .S2(n908), .D3(n899), .S3(n929), .Z(n2394) );
  HS65_LS_MX41X4 U12953 ( .D0(n838), .S0(n816), .D1(n840), .S1(n823), .D2(n833), .S2(n826), .D3(n817), .S3(n847), .Z(n1642) );
  HS65_LS_MX41X4 U12954 ( .D0(n879), .S0(n857), .D1(n881), .S1(n864), .D2(n874), .S2(n867), .D3(n858), .S3(n888), .Z(n1266) );
  HS65_LS_MX41X4 U12955 ( .D0(n797), .S0(n775), .D1(n799), .S1(n782), .D2(n792), .S2(n785), .D3(n776), .S3(n806), .Z(n2018) );
  HS65_LS_MX41X4 U12956 ( .D0(n167), .S0(n144), .D1(n155), .S1(n166), .D2(n156), .S2(n174), .D3(n165), .S3(n153), .Z(n4139) );
  HS65_LS_MX41X4 U12957 ( .D0(n200), .S0(n228), .D1(n212), .S1(n205), .D2(n217), .S2(n192), .D3(n222), .S3(n198), .Z(n3447) );
  HS65_LS_MX41X4 U12958 ( .D0(n332), .S0(n346), .D1(n327), .S1(n345), .D2(n318), .S2(n351), .D3(n358), .S3(n331), .Z(n8518) );
  HS65_LS_MX41X4 U12959 ( .D0(n807), .S0(n781), .D1(n798), .S1(n786), .D2(n778), .S2(n802), .D3(n772), .S3(n793), .Z(n2172) );
  HS65_LS_MX41X4 U12960 ( .D0(n889), .S0(n863), .D1(n880), .S1(n868), .D2(n860), .S2(n884), .D3(n854), .S3(n875), .Z(n1420) );
  HS65_LS_MX41X4 U12961 ( .D0(n848), .S0(n822), .D1(n839), .S1(n827), .D2(n819), .S2(n843), .D3(n813), .S3(n834), .Z(n1796) );
  HS65_LS_MX41X4 U12962 ( .D0(n930), .S0(n904), .D1(n921), .S1(n909), .D2(n901), .S2(n925), .D3(n895), .S3(n916), .Z(n2548) );
  HS65_LS_CB4I6X4 U12963 ( .A(n144), .B(n159), .C(n180), .D(n3564), .Z(n4096)
         );
  HS65_LS_MX41X4 U12964 ( .D0(n372), .S0(n391), .D1(n376), .S1(n387), .D2(n403), .S2(n373), .D3(n374), .S3(n397), .Z(n8226) );
  HS65_LS_CB4I6X4 U12965 ( .A(n572), .B(n573), .C(n536), .D(n6618), .Z(n6617)
         );
  HS65_LS_CB4I6X4 U12966 ( .A(n46), .B(n47), .C(n10), .D(n5025), .Z(n5024) );
  HS65_LS_CB4I6X4 U12967 ( .A(n76), .B(n73), .C(n68), .D(n6857), .Z(n6856) );
  HS65_LS_CB4I6X4 U12968 ( .A(n255), .B(n252), .C(n247), .D(n5265), .Z(n5264)
         );
  HS65_LS_CB4I6X4 U12969 ( .A(n474), .B(n471), .C(n466), .D(n5380), .Z(n5379)
         );
  HS65_LS_CB4I6X4 U12970 ( .A(n297), .B(n294), .C(n289), .D(n6972), .Z(n6971)
         );
  HS65_LS_CB4I6X4 U12971 ( .A(n710), .B(n711), .C(n675), .D(n5147), .Z(n5146)
         );
  HS65_LS_CB4I6X4 U12972 ( .A(n528), .B(n529), .C(n493), .D(n6739), .Z(n6738)
         );
  HS65_LS_MX41X4 U12973 ( .D0(n321), .S0(n341), .D1(n358), .S1(n330), .D2(n331), .S2(n354), .D3(n329), .S3(n350), .Z(n8874) );
  HS65_LS_MX41X4 U12974 ( .D0(n11), .S0(n29), .D1(n43), .S1(n26), .D2(n42), 
        .S2(n23), .D3(n24), .S3(n35), .Z(n5656) );
  HS65_LS_MX41X4 U12975 ( .D0(n537), .S0(n555), .D1(n569), .S1(n552), .D2(n568), .S2(n549), .D3(n550), .S3(n561), .Z(n7248) );
  HS65_LS_MX41X4 U12976 ( .D0(n165), .S0(n144), .D1(n156), .S1(n177), .D2(n176), .S2(n153), .D3(n154), .S3(n169), .Z(n4107) );
  HS65_LS_MX41X4 U12977 ( .D0(n479), .S0(n468), .D1(n485), .S1(n456), .D2(n489), .S2(n453), .D3(n484), .S3(n454), .Z(n5894) );
  HS65_LS_MX41X4 U12978 ( .D0(n260), .S0(n249), .D1(n266), .S1(n237), .D2(n270), .S2(n234), .D3(n265), .S3(n235), .Z(n5835) );
  HS65_LS_MX41X4 U12979 ( .D0(n693), .S0(n676), .D1(n707), .S1(n690), .D2(n706), .S2(n687), .D3(n699), .S3(n688), .Z(n5686) );
  HS65_LS_MX41X4 U12980 ( .D0(n302), .S0(n291), .D1(n308), .S1(n279), .D2(n312), .S2(n276), .D3(n307), .S3(n277), .Z(n7486) );
  HS65_LS_MX41X4 U12981 ( .D0(n81), .S0(n70), .D1(n87), .S1(n58), .D2(n91), 
        .S2(n55), .D3(n86), .S3(n56), .Z(n7427) );
  HS65_LS_MX41X4 U12982 ( .D0(n511), .S0(n494), .D1(n525), .S1(n508), .D2(n524), .S2(n505), .D3(n517), .S3(n506), .Z(n7278) );
  HS65_LS_MX41X4 U12983 ( .D0(n807), .S0(n772), .D1(n774), .S1(n802), .D2(n783), .S2(n793), .D3(n804), .S3(n773), .Z(n2212) );
  HS65_LS_MX41X4 U12984 ( .D0(n889), .S0(n854), .D1(n856), .S1(n884), .D2(n865), .S2(n875), .D3(n886), .S3(n855), .Z(n1460) );
  HS65_LS_MX41X4 U12985 ( .D0(n149), .S0(n176), .D1(n158), .S1(n180), .D2(n165), .S2(n150), .D3(n169), .S3(n157), .Z(n3558) );
  HS65_LS_MX41X4 U12986 ( .D0(n877), .S0(n865), .D1(n874), .S1(n853), .D2(n854), .S2(n887), .D3(n855), .S3(n885), .Z(n1276) );
  HS65_LS_MX41X4 U12987 ( .D0(n918), .S0(n906), .D1(n915), .S1(n894), .D2(n895), .S2(n928), .D3(n896), .S3(n926), .Z(n2404) );
  HS65_LS_MX41X4 U12988 ( .D0(n795), .S0(n783), .D1(n792), .S1(n771), .D2(n772), .S2(n805), .D3(n773), .S3(n803), .Z(n2028) );
  HS65_LS_MX41X4 U12989 ( .D0(n836), .S0(n824), .D1(n833), .S1(n812), .D2(n813), .S2(n846), .D3(n814), .S3(n844), .Z(n1652) );
  HS65_LS_MX41X4 U12990 ( .D0(n422), .S0(n445), .D1(n410), .S1(n432), .D2(n438), .S2(n421), .D3(n442), .S3(n412), .Z(n3793) );
  HS65_LS_MX41X4 U12991 ( .D0(n646), .S0(n669), .D1(n633), .S1(n656), .D2(n662), .S2(n645), .D3(n666), .S3(n635), .Z(n3676) );
  HS65_LS_MX41X4 U12992 ( .D0(n194), .S0(n223), .D1(n203), .S1(n226), .D2(n210), .S2(n195), .D3(n215), .S3(n202), .Z(n3432) );
  HS65_LS_IVX2 U12993 ( .A(n6939), .Z(n75) );
  HS65_LS_IVX2 U12994 ( .A(n6823), .Z(n516) );
  HS65_LS_IVX2 U12995 ( .A(n5231), .Z(n698) );
  HS65_LS_IVX2 U12996 ( .A(n5462), .Z(n473) );
  HS65_LS_IVX2 U12997 ( .A(n7054), .Z(n296) );
  HS65_LS_IVX2 U12998 ( .A(n5347), .Z(n254) );
  HS65_LS_AO212X4 U12999 ( .A(n420), .B(n3827), .C(n416), .D(n445), .E(n4346), 
        .Z(n4345) );
  HS65_LS_CB4I6X4 U13000 ( .A(n412), .B(n415), .C(n434), .D(n3899), .Z(n4346)
         );
  HS65_LS_AND3X4 U13001 ( .A(n4214), .B(n4215), .C(n4216), .Z(n4074) );
  HS65_LS_NOR4X4 U13002 ( .A(n3095), .B(n3108), .C(n3116), .D(n3455), .Z(n4215) );
  HS65_LS_NOR4ABX2 U13003 ( .A(n3466), .B(n2880), .C(n3478), .D(n3531), .Z(
        n4214) );
  HS65_LS_NOR4ABX2 U13004 ( .A(n4217), .B(n2952), .C(n3522), .D(n4218), .Z(
        n4216) );
  HS65_LS_AND3X4 U13005 ( .A(n4317), .B(n4318), .C(n4319), .Z(n3979) );
  HS65_LS_NOR4X4 U13006 ( .A(n3386), .B(n3397), .C(n3405), .D(n3815), .Z(n4318) );
  HS65_LS_NOR4ABX2 U13007 ( .A(n3826), .B(n3009), .C(n3837), .D(n3889), .Z(
        n4317) );
  HS65_LS_NOR4ABX2 U13008 ( .A(n4320), .B(n3195), .C(n3880), .D(n4321), .Z(
        n4319) );
  HS65_LS_AND3X4 U13009 ( .A(n4258), .B(n4259), .C(n4260), .Z(n3958) );
  HS65_LS_NOR4X4 U13010 ( .A(n3324), .B(n3335), .C(n3343), .D(n3698), .Z(n4259) );
  HS65_LS_NOR4ABX2 U13011 ( .A(n3761), .B(n3154), .C(n4261), .D(n4262), .Z(
        n4260) );
  HS65_LS_NOR4ABX2 U13012 ( .A(n3709), .B(n2991), .C(n3721), .D(n3772), .Z(
        n4258) );
  HS65_LS_OR3X4 U13013 ( .A(n1272), .B(n1273), .C(n1274), .Z(n1271) );
  HS65_LS_OR3X4 U13014 ( .A(n2024), .B(n2025), .C(n2026), .Z(n2023) );
  HS65_LS_OR3X4 U13015 ( .A(n2400), .B(n2401), .C(n2402), .Z(n2399) );
  HS65_LS_OR3X4 U13016 ( .A(n1648), .B(n1649), .C(n1650), .Z(n1647) );
  HS65_LS_OR3X4 U13017 ( .A(n3789), .B(n3790), .C(n3791), .Z(n3788) );
  HS65_LS_OA12X4 U13018 ( .A(n593), .B(n8400), .C(n623), .Z(n8398) );
  HS65_LS_OA12X4 U13019 ( .A(n106), .B(n8460), .C(n136), .Z(n8458) );
  HS65_LS_OA12X4 U13020 ( .A(n1604), .B(n845), .C(n824), .Z(n1781) );
  HS65_LS_OA12X4 U13021 ( .A(n2356), .B(n927), .C(n906), .Z(n2533) );
  HS65_LS_OA12X4 U13022 ( .A(n1980), .B(n804), .C(n783), .Z(n2157) );
  HS65_LS_OA12X4 U13023 ( .A(n1228), .B(n886), .C(n865), .Z(n1405) );
  HS65_LS_AO12X4 U13024 ( .A(n203), .B(n210), .C(n2936), .Z(n2935) );
  HS65_LS_AO12X4 U13025 ( .A(n410), .B(n438), .C(n3180), .Z(n3179) );
  HS65_LS_AO12X4 U13026 ( .A(n633), .B(n662), .C(n3139), .Z(n3138) );
  HS65_LS_AO12X4 U13027 ( .A(n158), .B(n165), .C(n3028), .Z(n3027) );
  HS65_LS_AO12X4 U13028 ( .A(n600), .B(n623), .C(n8142), .Z(n8141) );
  HS65_LS_AO12X4 U13029 ( .A(n113), .B(n136), .C(n8174), .Z(n8173) );
  HS65_LS_AO12X4 U13030 ( .A(n20), .B(n29), .C(n4552), .Z(n4551) );
  HS65_LS_AO12X4 U13031 ( .A(n546), .B(n555), .C(n6145), .Z(n6144) );
  HS65_LS_AO12X4 U13032 ( .A(n59), .B(n81), .C(n6330), .Z(n6329) );
  HS65_LS_AO12X4 U13033 ( .A(n457), .B(n479), .C(n4776), .Z(n4775) );
  HS65_LS_AO12X4 U13034 ( .A(n280), .B(n302), .C(n6369), .Z(n6368) );
  HS65_LS_AO12X4 U13035 ( .A(n238), .B(n260), .C(n4737), .Z(n4736) );
  HS65_LS_AO12X4 U13036 ( .A(n684), .B(n693), .C(n4629), .Z(n4628) );
  HS65_LS_AO12X4 U13037 ( .A(n502), .B(n511), .C(n6222), .Z(n6221) );
  HS65_LS_AO12X4 U13038 ( .A(n376), .B(n403), .C(n8011), .Z(n8010) );
  HS65_LS_AND3X4 U13039 ( .A(n6624), .B(n6160), .C(n6644), .Z(n7257) );
  HS65_LS_AND3X4 U13040 ( .A(n5031), .B(n4567), .C(n5051), .Z(n5665) );
  HS65_LS_OA12X4 U13041 ( .A(n7940), .B(n126), .C(n105), .Z(n7938) );
  HS65_LS_OA12X4 U13042 ( .A(n7841), .B(n613), .C(n592), .Z(n7839) );
  HS65_LS_OA12X4 U13043 ( .A(n8365), .B(n351), .C(n321), .Z(n8919) );
  HS65_LS_OA12X4 U13044 ( .A(n3268), .B(n172), .C(n144), .Z(n4128) );
  HS65_LS_NOR3AX2 U13045 ( .A(n6052), .B(n7448), .C(n7139), .Z(n7442) );
  HS65_LS_AO12X4 U13046 ( .A(n73), .B(n64), .C(n7135), .Z(n7448) );
  HS65_LS_NOR3AX2 U13047 ( .A(n7259), .B(n7260), .C(n7080), .Z(n7253) );
  HS65_LS_AO12X4 U13048 ( .A(n573), .B(n542), .C(n7266), .Z(n7260) );
  HS65_LS_NOR3AX2 U13049 ( .A(n5667), .B(n5668), .C(n5488), .Z(n5661) );
  HS65_LS_AO12X4 U13050 ( .A(n47), .B(n16), .C(n5674), .Z(n5668) );
  HS65_LS_NOR3AX2 U13051 ( .A(n4505), .B(n5915), .C(n5568), .Z(n5909) );
  HS65_LS_AO12X4 U13052 ( .A(n471), .B(n462), .C(n5564), .Z(n5915) );
  HS65_LS_NOR3AX2 U13053 ( .A(n6098), .B(n7507), .C(n7160), .Z(n7501) );
  HS65_LS_AO12X4 U13054 ( .A(n294), .B(n285), .C(n7156), .Z(n7507) );
  HS65_LS_NOR3AX2 U13055 ( .A(n4459), .B(n5856), .C(n5547), .Z(n5850) );
  HS65_LS_AO12X4 U13056 ( .A(n252), .B(n243), .C(n5543), .Z(n5856) );
  HS65_LS_NOR3AX2 U13057 ( .A(n5697), .B(n5698), .C(n5504), .Z(n5691) );
  HS65_LS_AO12X4 U13058 ( .A(n711), .B(n681), .C(n5704), .Z(n5698) );
  HS65_LS_NOR3AX2 U13059 ( .A(n7289), .B(n7290), .C(n7096), .Z(n7283) );
  HS65_LS_AO12X4 U13060 ( .A(n529), .B(n499), .C(n7296), .Z(n7290) );
  HS65_LS_OA12X4 U13061 ( .A(n3106), .B(n217), .C(n190), .Z(n4190) );
  HS65_LS_AO12X4 U13062 ( .A(n323), .B(n341), .C(n8053), .Z(n8052) );
  HS65_LS_OA12X4 U13063 ( .A(n1247), .B(n866), .C(n889), .Z(n1419) );
  HS65_LS_OA12X4 U13064 ( .A(n1999), .B(n784), .C(n807), .Z(n2171) );
  HS65_LS_OA12X4 U13065 ( .A(n1623), .B(n825), .C(n848), .Z(n1795) );
  HS65_LS_OA12X4 U13066 ( .A(n2375), .B(n907), .C(n930), .Z(n2547) );
  HS65_LS_OA12X4 U13067 ( .A(n4726), .B(n38), .C(n11), .Z(n5721) );
  HS65_LS_OA12X4 U13068 ( .A(n6319), .B(n564), .C(n537), .Z(n7313) );
  HS65_LS_OA12X4 U13069 ( .A(n4994), .B(n482), .C(n468), .Z(n5634) );
  HS65_LS_OA12X4 U13070 ( .A(n4940), .B(n263), .C(n249), .Z(n5607) );
  HS65_LS_OA12X4 U13071 ( .A(n6587), .B(n305), .C(n291), .Z(n7226) );
  HS65_LS_OA12X4 U13072 ( .A(n4866), .B(n702), .C(n676), .Z(n5783) );
  HS65_LS_OA12X4 U13073 ( .A(n6459), .B(n520), .C(n494), .Z(n7375) );
  HS65_LS_OA12X4 U13074 ( .A(n6533), .B(n84), .C(n70), .Z(n7199) );
  HS65_LS_OA12X4 U13075 ( .A(n8123), .B(n398), .C(n366), .Z(n8979) );
  HS65_LS_OA12X4 U13076 ( .A(n2922), .B(n157), .C(n170), .Z(n2921) );
  HS65_LS_OA12X4 U13077 ( .A(n7844), .B(n599), .C(n614), .Z(n7979) );
  HS65_LS_OA12X4 U13078 ( .A(n7883), .B(n112), .C(n127), .Z(n7992) );
  HS65_LS_OA12X4 U13079 ( .A(n6090), .B(n544), .C(n563), .Z(n6089) );
  HS65_LS_OA12X4 U13080 ( .A(n4497), .B(n18), .C(n37), .Z(n4496) );
  HS65_LS_OA12X4 U13081 ( .A(n1132), .B(n885), .C(n859), .Z(n1152) );
  HS65_LS_OA12X4 U13082 ( .A(n1884), .B(n803), .C(n777), .Z(n1904) );
  HS65_LS_OA12X4 U13083 ( .A(n3395), .B(n440), .C(n426), .Z(n4042) );
  HS65_LS_OA12X4 U13084 ( .A(n2852), .B(n412), .C(n441), .Z(n3001) );
  HS65_LS_OA12X4 U13085 ( .A(n4514), .B(n458), .C(n483), .Z(n4619) );
  HS65_LS_OA12X4 U13086 ( .A(n6107), .B(n281), .C(n306), .Z(n6212) );
  HS65_LS_OA12X4 U13087 ( .A(n6061), .B(n60), .C(n85), .Z(n6187) );
  HS65_LS_OA12X4 U13088 ( .A(n4468), .B(n239), .C(n264), .Z(n4594) );
  HS65_LS_OA12X4 U13089 ( .A(n2897), .B(n635), .C(n665), .Z(n2983) );
  HS65_LS_OA12X4 U13090 ( .A(n3333), .B(n664), .C(n650), .Z(n4018) );
  HS65_LS_OA12X4 U13091 ( .A(n7875), .B(n374), .C(n396), .Z(n7874) );
  HS65_LS_OA12X4 U13092 ( .A(n7958), .B(n324), .C(n353), .Z(n7957) );
  HS65_LS_IVX2 U13093 ( .A(n3553), .Z(n151) );
  HS65_LS_NOR3AX2 U13094 ( .A(n3554), .B(n3555), .C(n3556), .Z(n3553) );
  HS65_LS_IVX2 U13095 ( .A(n3671), .Z(n638) );
  HS65_LS_NOR3AX2 U13096 ( .A(n3672), .B(n3673), .C(n3674), .Z(n3671) );
  HS65_LS_IVX2 U13097 ( .A(n8769), .Z(n100) );
  HS65_LS_NOR3AX2 U13098 ( .A(n7921), .B(n8770), .C(n8771), .Z(n8769) );
  HS65_LS_IVX2 U13099 ( .A(n8681), .Z(n587) );
  HS65_LS_NOR3AX2 U13100 ( .A(n7822), .B(n8682), .C(n8683), .Z(n8681) );
  HS65_LS_IVX2 U13101 ( .A(n8514), .Z(n328) );
  HS65_LS_NOR3AX2 U13102 ( .A(n8515), .B(n8516), .C(n8517), .Z(n8514) );
  HS65_LS_IVX2 U13103 ( .A(n8155), .Z(n588) );
  HS65_LS_IVX2 U13104 ( .A(n8187), .Z(n101) );
  HS65_LS_OA12X4 U13105 ( .A(n350), .B(n8644), .C(n324), .Z(n8642) );
  HS65_LS_NAND3X2 U13106 ( .A(n9015), .B(n9016), .C(n9017), .Z(n7702) );
  HS65_LS_NOR4ABX2 U13107 ( .A(n8418), .B(n8740), .C(n8423), .D(n8408), .Z(
        n9016) );
  HS65_LS_NOR4ABX2 U13108 ( .A(n8695), .B(n7976), .C(n8729), .D(n8747), .Z(
        n9015) );
  HS65_LS_NOR4X4 U13109 ( .A(n8725), .B(n8156), .C(n9018), .D(n9019), .Z(n9017) );
  HS65_LS_NAND3X2 U13110 ( .A(n9073), .B(n9074), .C(n9075), .Z(n7740) );
  HS65_LS_NOR4ABX2 U13111 ( .A(n8478), .B(n8828), .C(n8483), .D(n8468), .Z(
        n9074) );
  HS65_LS_NOR4ABX2 U13112 ( .A(n8783), .B(n7989), .C(n8817), .D(n8835), .Z(
        n9073) );
  HS65_LS_NOR4X4 U13113 ( .A(n8813), .B(n8188), .C(n9076), .D(n9077), .Z(n9075) );
  HS65_LS_NAND3X2 U13114 ( .A(n7458), .B(n7459), .C(n7460), .Z(n7135) );
  HS65_LS_NOR4X4 U13115 ( .A(n6535), .B(n6924), .C(n6497), .D(n6523), .Z(n7459) );
  HS65_LS_NOR4ABX2 U13116 ( .A(n6866), .B(n6196), .C(n6913), .D(n6935), .Z(
        n7458) );
  HS65_LS_NOR4X4 U13117 ( .A(n6907), .B(n6350), .C(n7461), .D(n7462), .Z(n7460) );
  HS65_LS_NAND3X2 U13118 ( .A(n5925), .B(n5926), .C(n5927), .Z(n5564) );
  HS65_LS_NOR4X4 U13119 ( .A(n4996), .B(n5447), .C(n4958), .D(n4984), .Z(n5926) );
  HS65_LS_NOR4ABX2 U13120 ( .A(n5389), .B(n4615), .C(n5436), .D(n5458), .Z(
        n5925) );
  HS65_LS_NOR4X4 U13121 ( .A(n5430), .B(n4796), .C(n5928), .D(n5929), .Z(n5927) );
  HS65_LS_NAND3X2 U13122 ( .A(n7517), .B(n7518), .C(n7519), .Z(n7156) );
  HS65_LS_NOR4X4 U13123 ( .A(n6589), .B(n7039), .C(n6551), .D(n6577), .Z(n7518) );
  HS65_LS_NOR4ABX2 U13124 ( .A(n6981), .B(n6208), .C(n7028), .D(n7050), .Z(
        n7517) );
  HS65_LS_NOR4X4 U13125 ( .A(n7022), .B(n6389), .C(n7520), .D(n7521), .Z(n7519) );
  HS65_LS_NAND3X2 U13126 ( .A(n5866), .B(n5867), .C(n5868), .Z(n5543) );
  HS65_LS_NOR4X4 U13127 ( .A(n4942), .B(n5332), .C(n4904), .D(n4930), .Z(n5867) );
  HS65_LS_NOR4ABX2 U13128 ( .A(n5274), .B(n4603), .C(n5321), .D(n5343), .Z(
        n5866) );
  HS65_LS_NOR4X4 U13129 ( .A(n5315), .B(n4757), .C(n5869), .D(n5870), .Z(n5868) );
  HS65_LS_NAND3X2 U13130 ( .A(n5794), .B(n5795), .C(n5796), .Z(n5704) );
  HS65_LS_NOR4X4 U13131 ( .A(n4868), .B(n5216), .C(n4827), .D(n4854), .Z(n5795) );
  HS65_LS_NOR4ABX2 U13132 ( .A(n5157), .B(n4546), .C(n5205), .D(n5227), .Z(
        n5794) );
  HS65_LS_NOR4X4 U13133 ( .A(n5199), .B(n4650), .C(n5797), .D(n5798), .Z(n5796) );
  HS65_LS_NAND3X2 U13134 ( .A(n7386), .B(n7387), .C(n7388), .Z(n7296) );
  HS65_LS_NOR4X4 U13135 ( .A(n6461), .B(n6808), .C(n6420), .D(n6447), .Z(n7387) );
  HS65_LS_NOR4ABX2 U13136 ( .A(n6749), .B(n6139), .C(n6797), .D(n6819), .Z(
        n7386) );
  HS65_LS_NOR4X4 U13137 ( .A(n6791), .B(n6243), .C(n7389), .D(n7390), .Z(n7388) );
  HS65_LS_NAND3X2 U13138 ( .A(n7324), .B(n7325), .C(n7326), .Z(n7266) );
  HS65_LS_NOR4X4 U13139 ( .A(n6321), .B(n6687), .C(n6280), .D(n6307), .Z(n7325) );
  HS65_LS_NOR4ABX2 U13140 ( .A(n6677), .B(n6083), .C(n6629), .D(n6714), .Z(
        n7324) );
  HS65_LS_NOR4X4 U13141 ( .A(n6670), .B(n6166), .C(n7327), .D(n7328), .Z(n7326) );
  HS65_LS_NAND3X2 U13142 ( .A(n5732), .B(n5733), .C(n5734), .Z(n5674) );
  HS65_LS_NOR4X4 U13143 ( .A(n4728), .B(n5094), .C(n4687), .D(n4714), .Z(n5733) );
  HS65_LS_NOR4ABX2 U13144 ( .A(n5084), .B(n4490), .C(n5036), .D(n5121), .Z(
        n5732) );
  HS65_LS_NOR4X4 U13145 ( .A(n5077), .B(n4573), .C(n5735), .D(n5736), .Z(n5734) );
  HS65_LS_OA12X4 U13146 ( .A(n397), .B(n8506), .C(n374), .Z(n8674) );
  HS65_LS_NOR2X2 U13147 ( .A(n127), .B(n136), .Z(n7669) );
  HS65_LS_NOR2X2 U13148 ( .A(n191), .B(n204), .Z(n3126) );
  HS65_LS_NOR2X2 U13149 ( .A(n677), .B(n686), .Z(n4873) );
  HS65_LS_NOR2X2 U13150 ( .A(n495), .B(n504), .Z(n6466) );
  HS65_LS_OAI21X2 U13151 ( .A(n506), .B(n6426), .C(n524), .Z(n7099) );
  HS65_LS_OAI21X2 U13152 ( .A(n688), .B(n4833), .C(n706), .Z(n5507) );
  HS65_LS_OAI21X2 U13153 ( .A(n190), .B(n189), .C(n223), .Z(n2969) );
  HS65_LS_OAI21X2 U13154 ( .A(n357), .B(n353), .C(n337), .Z(n8887) );
  HS65_LS_OAI21X2 U13155 ( .A(n393), .B(n396), .C(n371), .Z(n9004) );
  HS65_LS_OAI21X2 U13156 ( .A(n566), .B(n563), .C(n542), .Z(n7120) );
  HS65_LS_OAI21X2 U13157 ( .A(n40), .B(n37), .C(n16), .Z(n5528) );
  HS65_LS_OAI21X2 U13158 ( .A(n126), .B(n136), .C(n112), .Z(n8446) );
  HS65_LS_OAI21X2 U13159 ( .A(n357), .B(n344), .C(n336), .Z(n8327) );
  HS65_LS_OAI21X2 U13160 ( .A(n662), .B(n670), .C(n648), .Z(n2988) );
  HS65_LS_OAI21X2 U13161 ( .A(n341), .B(n356), .C(n322), .Z(n7962) );
  HS65_LS_OAI21X2 U13162 ( .A(n702), .B(n693), .C(n683), .Z(n4878) );
  HS65_LS_OAI21X2 U13163 ( .A(n217), .B(n210), .C(n202), .Z(n3131) );
  HS65_LS_OAI21X2 U13164 ( .A(n351), .B(n341), .C(n324), .Z(n8330) );
  HS65_LS_OAI21X2 U13165 ( .A(n83), .B(n74), .C(n69), .Z(n6363) );
  HS65_LS_OAI21X2 U13166 ( .A(n481), .B(n472), .C(n467), .Z(n4809) );
  HS65_LS_OAI21X2 U13167 ( .A(n304), .B(n295), .C(n290), .Z(n6402) );
  HS65_LS_OAI21X2 U13168 ( .A(n262), .B(n253), .C(n248), .Z(n4770) );
  HS65_LS_OAI21X2 U13169 ( .A(n700), .B(n712), .C(n677), .Z(n4663) );
  HS65_LS_OAI21X2 U13170 ( .A(n518), .B(n530), .C(n495), .Z(n6256) );
  HS65_LS_OAI21X2 U13171 ( .A(n615), .B(n609), .C(n589), .Z(n8168) );
  HS65_LS_OAI21X2 U13172 ( .A(n128), .B(n122), .C(n102), .Z(n8200) );
  HS65_LS_OAI21X2 U13173 ( .A(n70), .B(n68), .C(n91), .Z(n6362) );
  HS65_LS_OAI21X2 U13174 ( .A(n291), .B(n289), .C(n312), .Z(n6401) );
  HS65_LS_OAI21X2 U13175 ( .A(n249), .B(n247), .C(n270), .Z(n4769) );
  HS65_LS_OAI21X2 U13176 ( .A(n676), .B(n675), .C(n706), .Z(n4662) );
  HS65_LS_OAI21X2 U13177 ( .A(n494), .B(n493), .C(n524), .Z(n6255) );
  HS65_LS_OAI21X2 U13178 ( .A(n366), .B(n369), .C(n391), .Z(n8007) );
  HS65_LS_OAI21X2 U13179 ( .A(n321), .B(n322), .C(n354), .Z(n8049) );
  HS65_LS_OAI21X2 U13180 ( .A(n426), .B(n424), .C(n445), .Z(n3212) );
  HS65_LS_OAI21X2 U13181 ( .A(n592), .B(n591), .C(n618), .Z(n8167) );
  HS65_LS_OAI21X2 U13182 ( .A(n105), .B(n104), .C(n131), .Z(n8199) );
  HS65_LS_NOR2X2 U13183 ( .A(n352), .B(n343), .Z(n8325) );
  HS65_LS_BFX2 U13184 ( .A(n9148), .Z(n9142) );
  HS65_LS_IVX2 U13185 ( .A(n3467), .Z(n211) );
  HS65_LS_IVX2 U13186 ( .A(n3292), .Z(n146) );
  HS65_LS_IVX2 U13187 ( .A(n8249), .Z(n389) );
  HS65_LS_IVX2 U13188 ( .A(n8553), .Z(n342) );
  HS65_LS_IVX2 U13190 ( .A(n5086), .Z(n30) );
  HS65_LS_IVX2 U13191 ( .A(n6679), .Z(n556) );
  HS65_LS_IVX2 U13192 ( .A(n6800), .Z(n512) );
  HS65_LS_IVX2 U13193 ( .A(n5208), .Z(n694) );
  HS65_LS_IVX2 U13194 ( .A(n7758), .Z(n368) );
  HS65_LS_IVX2 U13195 ( .A(n7775), .Z(n320) );
  HS65_LS_IVX2 U13196 ( .A(n4671), .Z(n13) );
  HS65_LS_IVX2 U13197 ( .A(n6264), .Z(n539) );
  HS65_LS_IVX2 U13198 ( .A(n7684), .Z(n590) );
  HS65_LS_IVX2 U13199 ( .A(n7722), .Z(n103) );
  HS65_LS_OA12X4 U13202 ( .A(n3247), .B(n154), .C(n176), .Z(n3920) );
  HS65_LS_OA12X4 U13203 ( .A(n4537), .B(n683), .C(n701), .Z(n4536) );
  HS65_LS_OA12X4 U13204 ( .A(n6130), .B(n501), .C(n519), .Z(n6129) );
  HS65_LS_OA12X4 U13205 ( .A(n2872), .B(n202), .C(n216), .Z(n2871) );
  HS65_LS_NAND2X2 U13207 ( .A(n2592), .B(n2593), .Z(n2264) );
  HS65_LS_NAND2X2 U13208 ( .A(n2216), .B(n2217), .Z(n1888) );
  HS65_LS_NAND2X2 U13209 ( .A(n1840), .B(n1841), .Z(n1512) );
  HS65_LS_NAND2X2 U13210 ( .A(n1464), .B(n1465), .Z(n1136) );
  HS65_LS_NAND2X2 U13211 ( .A(n4222), .B(n4212), .Z(n2878) );
  HS65_LS_NAND2X2 U13212 ( .A(n8998), .B(n8999), .Z(n7862) );
  HS65_LS_NAND4ABX3 U13213 ( .A(n8443), .B(n8444), .C(n8445), .D(n8446), .Z(
        n8439) );
  HS65_LS_OAI212X3 U13214 ( .A(n8441), .B(n7660), .C(n103), .D(n7667), .E(
        n8442), .Z(n8440) );
  HS65_LS_AOI212X2 U13215 ( .A(n113), .B(n8448), .C(n110), .D(n122), .E(n8449), 
        .Z(n8438) );
  HS65_LS_NOR4ABX2 U13216 ( .A(n8035), .B(n8036), .C(n8037), .D(n8038), .Z(
        n3013) );
  HS65_LS_NAND4ABX3 U13217 ( .A(n8047), .B(n8048), .C(n8049), .D(n8050), .Z(
        n8037) );
  HS65_LS_OAI212X3 U13218 ( .A(n8039), .B(n8040), .C(n8041), .D(n7964), .E(
        n8042), .Z(n8038) );
  HS65_LS_AOI212X2 U13219 ( .A(n350), .B(n322), .C(n335), .D(n345), .E(n8052), 
        .Z(n8036) );
  HS65_LS_NOR4ABX2 U13220 ( .A(n7967), .B(n7968), .C(n7969), .D(n7970), .Z(
        n2791) );
  HS65_LS_CBI4I1X3 U13221 ( .A(n7697), .B(n7817), .C(n7641), .D(n7976), .Z(
        n7969) );
  HS65_LS_CBI4I6X2 U13222 ( .A(n593), .B(n7709), .C(n624), .D(n7977), .Z(n7968) );
  HS65_LS_AOI212X2 U13223 ( .A(n608), .B(n586), .C(n596), .D(n618), .E(n7979), 
        .Z(n7967) );
  HS65_LS_NOR4ABX2 U13224 ( .A(n5648), .B(n5649), .C(n5650), .D(n5651), .Z(
        n2777) );
  HS65_LS_MX41X4 U13225 ( .D0(n38), .S0(n16), .D1(n48), .S1(n23), .D2(n24), 
        .S2(n37), .D3(n17), .S3(n4571), .Z(n5651) );
  HS65_LS_MX41X4 U13226 ( .D0(n36), .S0(n4491), .D1(n10), .S1(n32), .D2(n14), 
        .S2(n47), .D3(n33), .S3(n20), .Z(n5650) );
  HS65_LS_NOR4ABX2 U13227 ( .A(n5053), .B(n5652), .C(n5033), .D(n4564), .Z(
        n5649) );
  HS65_LS_NOR4ABX2 U13228 ( .A(n7240), .B(n7241), .C(n7242), .D(n7243), .Z(
        n2769) );
  HS65_LS_MX41X4 U13229 ( .D0(n564), .S0(n542), .D1(n574), .S1(n549), .D2(n550), .S2(n563), .D3(n543), .S3(n6164), .Z(n7243) );
  HS65_LS_MX41X4 U13230 ( .D0(n562), .S0(n6084), .D1(n536), .S1(n558), .D2(
        n540), .S2(n573), .D3(n559), .S3(n546), .Z(n7242) );
  HS65_LS_NOR4ABX2 U13231 ( .A(n6646), .B(n7244), .C(n6626), .D(n6157), .Z(
        n7241) );
  HS65_LS_NAND4ABX3 U13232 ( .A(n7887), .B(n7888), .C(n7889), .D(n7890), .Z(
        n7878) );
  HS65_LS_OAI212X3 U13233 ( .A(n7725), .B(n7880), .C(n7660), .D(n7881), .E(
        n7882), .Z(n7879) );
  HS65_LS_AOI212X2 U13234 ( .A(n106), .B(n127), .C(n119), .D(n114), .E(n7892), 
        .Z(n7877) );
  HS65_LS_NOR4ABX2 U13235 ( .A(n4664), .B(n4665), .C(n4666), .D(n4667), .Z(
        n2781) );
  HS65_LS_NAND4ABX3 U13236 ( .A(n4672), .B(n4673), .C(n4674), .D(n4675), .Z(
        n4666) );
  HS65_LS_OAI212X3 U13237 ( .A(n4668), .B(n4560), .C(n13), .D(n4669), .E(n4670), .Z(n4667) );
  HS65_LS_AOI212X2 U13238 ( .A(n20), .B(n4678), .C(n48), .D(n23), .E(n4679), 
        .Z(n4665) );
  HS65_LS_CBI4I1X3 U13239 ( .A(n2966), .B(n3100), .C(n2874), .D(n3509), .Z(
        n3902) );
  HS65_LS_AOI212X2 U13240 ( .A(n217), .B(n202), .C(n203), .D(n3911), .E(n3912), 
        .Z(n3900) );
  HS65_LS_CBI4I1X3 U13241 ( .A(n211), .B(n3102), .C(n2877), .D(n3904), .Z(
        n3903) );
  HS65_LS_CBI4I6X2 U13242 ( .A(n455), .B(n4616), .C(n480), .D(n4617), .Z(n4605) );
  HS65_LS_CBI4I1X3 U13243 ( .A(n4613), .B(n4510), .C(n4614), .D(n4615), .Z(
        n4606) );
  HS65_LS_AOI212X2 U13244 ( .A(n474), .B(n463), .C(n489), .D(n456), .E(n4619), 
        .Z(n4604) );
  HS65_LS_CBI4I6X2 U13245 ( .A(n278), .B(n6209), .C(n303), .D(n6210), .Z(n6198) );
  HS65_LS_CBI4I1X3 U13246 ( .A(n6206), .B(n6103), .C(n6207), .D(n6208), .Z(
        n6199) );
  HS65_LS_AOI212X2 U13247 ( .A(n297), .B(n286), .C(n312), .D(n279), .E(n6212), 
        .Z(n6197) );
  HS65_LS_CBI4I1X3 U13248 ( .A(n7735), .B(n7880), .C(n7669), .D(n7989), .Z(
        n7982) );
  HS65_LS_CBI4I6X2 U13249 ( .A(n106), .B(n7747), .C(n137), .D(n7990), .Z(n7981) );
  HS65_LS_AOI212X2 U13250 ( .A(n121), .B(n99), .C(n109), .D(n131), .E(n7992), 
        .Z(n7980) );
  HS65_LS_NOR4ABX2 U13251 ( .A(n6257), .B(n6258), .C(n6259), .D(n6260), .Z(
        n2773) );
  HS65_LS_NAND4ABX3 U13252 ( .A(n6265), .B(n6266), .C(n6267), .D(n6268), .Z(
        n6259) );
  HS65_LS_OAI212X3 U13253 ( .A(n6261), .B(n6153), .C(n539), .D(n6262), .E(
        n6263), .Z(n6260) );
  HS65_LS_AOI212X2 U13254 ( .A(n546), .B(n6271), .C(n574), .D(n549), .E(n6272), 
        .Z(n6258) );
  HS65_LS_NOR4ABX2 U13255 ( .A(n7993), .B(n7994), .C(n7995), .D(n7996), .Z(
        n2766) );
  HS65_LS_NAND4ABX3 U13256 ( .A(n8005), .B(n8006), .C(n8007), .D(n8008), .Z(
        n7995) );
  HS65_LS_OAI212X3 U13257 ( .A(n7997), .B(n7998), .C(n7999), .D(n7862), .E(
        n8000), .Z(n7996) );
  HS65_LS_AOI212X2 U13258 ( .A(n397), .B(n369), .C(n370), .D(n404), .E(n8010), 
        .Z(n7994) );
  HS65_LS_NOR4ABX2 U13259 ( .A(n6071), .B(n6072), .C(n6073), .D(n6074), .Z(
        n2775) );
  HS65_LS_CBI4I6X2 U13260 ( .A(n551), .B(n6084), .C(n557), .D(n6085), .Z(n6072) );
  HS65_LS_CBI4I1X3 U13261 ( .A(n6080), .B(n6081), .C(n6082), .D(n6083), .Z(
        n6073) );
  HS65_LS_AOI212X2 U13262 ( .A(n543), .B(n572), .C(n568), .D(n552), .E(n6089), 
        .Z(n6071) );
  HS65_LS_NOR4ABX2 U13263 ( .A(n8321), .B(n8322), .C(n8323), .D(n8324), .Z(
        n3012) );
  HS65_LS_NAND4ABX3 U13264 ( .A(n8328), .B(n8329), .C(n8330), .D(n8331), .Z(
        n8323) );
  HS65_LS_OAI212X3 U13265 ( .A(n8325), .B(n7955), .C(n320), .D(n8326), .E(
        n8327), .Z(n8324) );
  HS65_LS_AOI212X2 U13266 ( .A(n323), .B(n8333), .C(n331), .D(n346), .E(n8334), 
        .Z(n8322) );
  HS65_LS_NOR4ABX2 U13267 ( .A(n4478), .B(n4479), .C(n4480), .D(n4481), .Z(
        n2783) );
  HS65_LS_CBI4I6X2 U13268 ( .A(n25), .B(n4491), .C(n31), .D(n4492), .Z(n4479)
         );
  HS65_LS_CBI4I1X3 U13269 ( .A(n4487), .B(n4488), .C(n4489), .D(n4490), .Z(
        n4480) );
  HS65_LS_AOI212X2 U13270 ( .A(n17), .B(n46), .C(n42), .D(n26), .E(n4496), .Z(
        n4478) );
  HS65_LS_NOR4ABX2 U13271 ( .A(n7853), .B(n7854), .C(n7855), .D(n7856), .Z(
        n2767) );
  HS65_LS_CBI4I1X3 U13272 ( .A(n7857), .B(n7858), .C(n7859), .D(n7860), .Z(
        n7856) );
  HS65_LS_CBI4I1X3 U13273 ( .A(n7861), .B(n7862), .C(n7863), .D(n7864), .Z(
        n7855) );
  HS65_LS_AOI212X2 U13274 ( .A(n387), .B(n373), .C(n379), .D(n391), .E(n7874), 
        .Z(n7853) );
  HS65_LS_NOR4ABX2 U13275 ( .A(n8883), .B(n8884), .C(n8885), .D(n8886), .Z(
        n2630) );
  HS65_LS_CB4I6X4 U13276 ( .A(n344), .B(n343), .C(n324), .D(n8591), .Z(n8885)
         );
  HS65_LS_CBI4I1X3 U13277 ( .A(n7965), .B(n7954), .C(n7778), .D(n8887), .Z(
        n8886) );
  HS65_LS_AOI222X2 U13278 ( .A(n334), .B(n350), .C(n323), .D(n8943), .E(n341), 
        .F(n329), .Z(n8883) );
  HS65_LS_IVX2 U13279 ( .A(n4680), .Z(n12) );
  HS65_LS_IVX2 U13280 ( .A(n6273), .Z(n538) );
  HS65_LS_IVX2 U13281 ( .A(n3067), .Z(n145) );
  HS65_LS_NOR4ABX2 U13282 ( .A(n6475), .B(n6476), .C(n6477), .D(n6478), .Z(
        n2797) );
  HS65_LS_NAND4ABX3 U13283 ( .A(n6483), .B(n6484), .C(n6485), .D(n6486), .Z(
        n6477) );
  HS65_LS_OAI212X3 U13284 ( .A(n6479), .B(n6058), .C(n6480), .D(n6481), .E(
        n6482), .Z(n6478) );
  HS65_LS_AOI212X2 U13285 ( .A(n59), .B(n6489), .C(n74), .D(n55), .E(n6490), 
        .Z(n6476) );
  HS65_LS_NOR4ABX2 U13286 ( .A(n4882), .B(n4883), .C(n4884), .D(n4885), .Z(
        n2805) );
  HS65_LS_NAND4ABX3 U13287 ( .A(n4890), .B(n4891), .C(n4892), .D(n4893), .Z(
        n4884) );
  HS65_LS_OAI212X3 U13288 ( .A(n4886), .B(n4465), .C(n4887), .D(n4888), .E(
        n4889), .Z(n4885) );
  HS65_LS_AOI212X2 U13289 ( .A(n238), .B(n4896), .C(n253), .D(n234), .E(n4897), 
        .Z(n4883) );
  HS65_LS_IVX2 U13290 ( .A(n7760), .Z(n367) );
  HS65_LS_IVX2 U13291 ( .A(n7777), .Z(n319) );
  HS65_LS_NAND4ABX3 U13292 ( .A(n5767), .B(n5768), .C(n5769), .D(n5770), .Z(
        n3544) );
  HS65_LS_NAND4ABX3 U13293 ( .A(n5183), .B(n5233), .C(n5827), .D(n5828), .Z(
        n5767) );
  HS65_LS_OAI212X3 U13294 ( .A(n4862), .B(n4544), .C(n4636), .D(n4860), .E(
        n5825), .Z(n5768) );
  HS65_LS_AOI212X2 U13295 ( .A(n689), .B(n701), .C(n685), .D(n709), .E(n5771), 
        .Z(n5770) );
  HS65_LS_NAND4ABX3 U13296 ( .A(n7359), .B(n7360), .C(n7361), .D(n7362), .Z(
        n3219) );
  HS65_LS_NAND4ABX3 U13297 ( .A(n6775), .B(n6825), .C(n7419), .D(n7420), .Z(
        n7359) );
  HS65_LS_OAI212X3 U13298 ( .A(n6455), .B(n6137), .C(n6229), .D(n6453), .E(
        n7417), .Z(n7360) );
  HS65_LS_AOI212X2 U13299 ( .A(n507), .B(n519), .C(n503), .D(n527), .E(n7363), 
        .Z(n7362) );
  HS65_LS_NAND4ABX3 U13300 ( .A(n4452), .B(n4453), .C(n4454), .D(n4455), .Z(
        n2808) );
  HS65_LS_NAND4ABX3 U13301 ( .A(n4473), .B(n4474), .C(n4475), .D(n4476), .Z(
        n4452) );
  HS65_LS_OAI212X3 U13302 ( .A(n4463), .B(n4464), .C(n4465), .D(n4466), .E(
        n4467), .Z(n4453) );
  HS65_LS_AOI212X2 U13303 ( .A(n236), .B(n264), .C(n240), .D(n256), .E(n4456), 
        .Z(n4455) );
  HS65_LS_NAND4ABX3 U13304 ( .A(n6045), .B(n6046), .C(n6047), .D(n6048), .Z(
        n2800) );
  HS65_LS_NAND4ABX3 U13305 ( .A(n6066), .B(n6067), .C(n6068), .D(n6069), .Z(
        n6045) );
  HS65_LS_OAI212X3 U13306 ( .A(n6056), .B(n6057), .C(n6058), .D(n6059), .E(
        n6060), .Z(n6046) );
  HS65_LS_AOI212X2 U13307 ( .A(n57), .B(n85), .C(n61), .D(n77), .E(n6049), .Z(
        n6048) );
  HS65_LS_NAND4ABX3 U13308 ( .A(n7088), .B(n7089), .C(n7090), .D(n7091), .Z(
        n3018) );
  HS65_LS_AOI212X2 U13309 ( .A(n501), .B(n520), .C(n502), .D(n7097), .E(n7098), 
        .Z(n7090) );
  HS65_LS_CBI4I1X3 U13310 ( .A(n6252), .B(n6453), .C(n6452), .D(n6773), .Z(
        n7088) );
  HS65_LS_CBI4I1X3 U13311 ( .A(n512), .B(n6455), .C(n6136), .D(n7099), .Z(
        n7089) );
  HS65_LS_NAND4ABX3 U13312 ( .A(n5496), .B(n5497), .C(n5498), .D(n5499), .Z(
        n3222) );
  HS65_LS_AOI212X2 U13313 ( .A(n683), .B(n702), .C(n684), .D(n5505), .E(n5506), 
        .Z(n5498) );
  HS65_LS_CBI4I1X3 U13314 ( .A(n4659), .B(n4860), .C(n4859), .D(n5181), .Z(
        n5496) );
  HS65_LS_CBI4I1X3 U13315 ( .A(n694), .B(n4862), .C(n4543), .D(n5507), .Z(
        n5497) );
  HS65_LS_NAND4ABX3 U13316 ( .A(n8855), .B(n8856), .C(n8857), .D(n8858), .Z(
        n3010) );
  HS65_LS_AOI212X2 U13317 ( .A(n324), .B(n351), .C(n323), .D(n8644), .E(n8880), 
        .Z(n8857) );
  HS65_LS_CB4I6X4 U13318 ( .A(n344), .B(n350), .C(n332), .D(n8589), .Z(n8855)
         );
  HS65_LS_CBI4I1X3 U13319 ( .A(n342), .B(n7779), .C(n7963), .D(n8882), .Z(
        n8856) );
  HS65_LS_NAND4ABX3 U13320 ( .A(n7788), .B(n7789), .C(n7790), .D(n7791), .Z(
        n2792) );
  HS65_LS_OAI212X3 U13321 ( .A(n7687), .B(n7817), .C(n7632), .D(n7842), .E(
        n7843), .Z(n7789) );
  HS65_LS_NAND4ABX3 U13322 ( .A(n7848), .B(n7849), .C(n7850), .D(n7851), .Z(
        n7788) );
  HS65_LS_AOI212X2 U13323 ( .A(n593), .B(n614), .C(n606), .D(n601), .E(n7792), 
        .Z(n7791) );
  HS65_LS_NAND4ABX3 U13324 ( .A(n4112), .B(n4113), .C(n4114), .D(n4115), .Z(
        n2691) );
  HS65_LS_NAND4ABX3 U13325 ( .A(n3645), .B(n3578), .C(n4172), .D(n4173), .Z(
        n4112) );
  HS65_LS_OAI212X3 U13326 ( .A(n3264), .B(n2928), .C(n3042), .D(n3262), .E(
        n4170), .Z(n4113) );
  HS65_LS_AOI212X2 U13327 ( .A(n170), .B(n155), .C(n160), .D(n179), .E(n4116), 
        .Z(n4115) );
  HS65_LS_NAND4ABX3 U13328 ( .A(n5678), .B(n5679), .C(n5680), .D(n5681), .Z(
        n3220) );
  HS65_LS_MX41X4 U13329 ( .D0(n702), .S0(n681), .D1(n712), .S1(n687), .D2(n688), .S2(n701), .D3(n682), .S3(n4648), .Z(n5679) );
  HS65_LS_MX41X4 U13330 ( .D0(n700), .S0(n4531), .D1(n675), .S1(n696), .D2(
        n679), .S2(n711), .D3(n697), .S3(n684), .Z(n5678) );
  HS65_LS_NOR4ABX2 U13331 ( .A(n5173), .B(n5154), .C(n5682), .D(n4641), .Z(
        n5681) );
  HS65_LS_NAND4ABX3 U13332 ( .A(n7270), .B(n7271), .C(n7272), .D(n7273), .Z(
        n3016) );
  HS65_LS_MX41X4 U13333 ( .D0(n520), .S0(n499), .D1(n530), .S1(n505), .D2(n506), .S2(n519), .D3(n500), .S3(n6241), .Z(n7271) );
  HS65_LS_MX41X4 U13334 ( .D0(n518), .S0(n6124), .D1(n493), .S1(n514), .D2(
        n497), .S2(n529), .D3(n515), .S3(n502), .Z(n7270) );
  HS65_LS_NOR4ABX2 U13335 ( .A(n6765), .B(n6746), .C(n7274), .D(n6234), .Z(
        n7273) );
  HS65_LS_NAND4ABX3 U13336 ( .A(n4174), .B(n4175), .C(n4176), .D(n4177), .Z(
        n2732) );
  HS65_LS_NAND4ABX3 U13337 ( .A(n3498), .B(n3532), .C(n4234), .D(n4235), .Z(
        n4174) );
  HS65_LS_OAI212X3 U13338 ( .A(n3102), .B(n2878), .C(n3100), .D(n2943), .E(
        n4232), .Z(n4175) );
  HS65_LS_AOI212X2 U13339 ( .A(n200), .B(n216), .C(n205), .D(n225), .E(n4178), 
        .Z(n4177) );
  HS65_LS_NAND4ABX3 U13340 ( .A(n7676), .B(n7677), .C(n7678), .D(n7679), .Z(
        n2785) );
  HS65_LS_NOR4ABX2 U13341 ( .A(n7680), .B(n7681), .C(n7682), .D(n7683), .Z(
        n7679) );
  HS65_LS_MX41X4 U13342 ( .D0(n613), .S0(n583), .D1(n597), .S1(n609), .D2(n594), .S2(n614), .D3(n586), .S3(n7710), .Z(n7677) );
  HS65_LS_MX41X4 U13343 ( .D0(n615), .S0(n7709), .D1(n591), .S1(n625), .D2(
        n585), .S2(n611), .D3(n622), .S3(n600), .Z(n7676) );
  HS65_LS_NAND4ABX3 U13344 ( .A(n8645), .B(n8646), .C(n8647), .D(n8648), .Z(
        n2768) );
  HS65_LS_OAI212X3 U13345 ( .A(n7862), .B(n7762), .C(n8119), .D(n7872), .E(
        n8672), .Z(n8646) );
  HS65_LS_NAND4ABX3 U13346 ( .A(n8674), .B(n8311), .C(n8275), .D(n8675), .Z(
        n8645) );
  HS65_LS_AOI212X2 U13347 ( .A(n381), .B(n396), .C(n375), .D(n388), .E(n8649), 
        .Z(n8648) );
  HS65_LS_IVX2 U13348 ( .A(n2328), .Z(n924) );
  HS65_LS_IVX2 U13349 ( .A(n1576), .Z(n842) );
  HS65_LS_IVX2 U13350 ( .A(n1952), .Z(n801) );
  HS65_LS_IVX2 U13351 ( .A(n1200), .Z(n883) );
  HS65_LS_NAND4ABX3 U13352 ( .A(n2881), .B(n2882), .C(n2883), .D(n2884), .Z(
        n2639) );
  HS65_LS_NAND4ABX3 U13353 ( .A(n2902), .B(n2903), .C(n2904), .D(n2905), .Z(
        n2881) );
  HS65_LS_OAI212X3 U13354 ( .A(n2892), .B(n2893), .C(n2894), .D(n2895), .E(
        n2896), .Z(n2882) );
  HS65_LS_AOI212X2 U13355 ( .A(n641), .B(n665), .C(n634), .D(n658), .E(n2885), 
        .Z(n2884) );
  HS65_LS_IVX2 U13356 ( .A(n6080), .Z(n548) );
  HS65_LS_IVX2 U13357 ( .A(n4487), .Z(n22) );
  HS65_LS_NAND4ABX3 U13358 ( .A(n4624), .B(n4625), .C(n4626), .D(n4627), .Z(
        n3225) );
  HS65_LS_NAND4ABX3 U13359 ( .A(n4660), .B(n4661), .C(n4662), .D(n4663), .Z(
        n4624) );
  HS65_LS_OAI212X3 U13360 ( .A(n4652), .B(n4653), .C(n4544), .D(n4654), .E(
        n4655), .Z(n4625) );
  HS65_LS_AOI212X2 U13361 ( .A(n675), .B(n699), .C(n695), .D(n679), .E(n4628), 
        .Z(n4627) );
  HS65_LS_NAND4ABX3 U13362 ( .A(n6217), .B(n6218), .C(n6219), .D(n6220), .Z(
        n3217) );
  HS65_LS_NAND4ABX3 U13363 ( .A(n6253), .B(n6254), .C(n6255), .D(n6256), .Z(
        n6217) );
  HS65_LS_OAI212X3 U13364 ( .A(n6245), .B(n6246), .C(n6137), .D(n6247), .E(
        n6248), .Z(n6218) );
  HS65_LS_AOI212X2 U13365 ( .A(n493), .B(n517), .C(n513), .D(n497), .E(n6221), 
        .Z(n6220) );
  HS65_LS_NAND4ABX3 U13366 ( .A(n7944), .B(n7945), .C(n7946), .D(n7947), .Z(
        n3014) );
  HS65_LS_CBI4I1X3 U13367 ( .A(n7959), .B(n7960), .C(n7961), .D(n7962), .Z(
        n7945) );
  HS65_LS_CBI4I1X3 U13368 ( .A(n7963), .B(n7964), .C(n7965), .D(n7966), .Z(
        n7944) );
  HS65_LS_AOI212X2 U13369 ( .A(n347), .B(n336), .C(n330), .D(n354), .E(n7957), 
        .Z(n7946) );
  HS65_LS_IVX2 U13370 ( .A(n7871), .Z(n386) );
  HS65_LS_NAND4ABX3 U13371 ( .A(n6539), .B(n6540), .C(n6541), .D(n6542), .Z(
        n2821) );
  HS65_LS_NAND4ABX3 U13372 ( .A(n6597), .B(n6598), .C(n6599), .D(n6600), .Z(
        n6539) );
  HS65_LS_OAI212X3 U13373 ( .A(n6593), .B(n6104), .C(n6594), .D(n6595), .E(
        n6596), .Z(n6540) );
  HS65_LS_AOI212X2 U13374 ( .A(n280), .B(n6543), .C(n295), .D(n276), .E(n6544), 
        .Z(n6542) );
  HS65_LS_NAND4ABX3 U13375 ( .A(n4946), .B(n4947), .C(n4948), .D(n4949), .Z(
        n2829) );
  HS65_LS_NAND4ABX3 U13376 ( .A(n5004), .B(n5005), .C(n5006), .D(n5007), .Z(
        n4946) );
  HS65_LS_OAI212X3 U13377 ( .A(n5000), .B(n4511), .C(n5001), .D(n5002), .E(
        n5003), .Z(n4947) );
  HS65_LS_AOI212X2 U13378 ( .A(n457), .B(n4950), .C(n472), .D(n453), .E(n4951), 
        .Z(n4949) );
  HS65_LS_NAND4ABX3 U13379 ( .A(n3175), .B(n3176), .C(n3177), .D(n3178), .Z(
        n2701) );
  HS65_LS_NAND4ABX3 U13380 ( .A(n3210), .B(n3211), .C(n3212), .D(n3213), .Z(
        n3175) );
  HS65_LS_OAI212X3 U13381 ( .A(n3202), .B(n3203), .C(n3204), .D(n2848), .E(
        n3205), .Z(n3176) );
  HS65_LS_AOI212X2 U13382 ( .A(n424), .B(n442), .C(n419), .D(n437), .E(n3179), 
        .Z(n3178) );
  HS65_LS_NAND4ABX3 U13383 ( .A(n3023), .B(n3024), .C(n3025), .D(n3026), .Z(
        n2646) );
  HS65_LS_NAND4ABX3 U13384 ( .A(n3059), .B(n3060), .C(n3061), .D(n3062), .Z(
        n3023) );
  HS65_LS_OAI212X3 U13385 ( .A(n3051), .B(n3052), .C(n3053), .D(n2928), .E(
        n3054), .Z(n3024) );
  HS65_LS_AOI212X2 U13386 ( .A(n143), .B(n169), .C(n148), .D(n166), .E(n3027), 
        .Z(n3026) );
  HS65_LS_IVX2 U13387 ( .A(n3044), .Z(n181) );
  HS65_LS_NAND4ABX3 U13388 ( .A(n5621), .B(n5622), .C(n5623), .D(n5624), .Z(
        n2826) );
  HS65_LS_CB4I6X4 U13389 ( .A(n478), .B(n477), .C(n458), .D(n5416), .Z(n5621)
         );
  HS65_LS_CBI4I1X3 U13390 ( .A(n4614), .B(n5565), .C(n5645), .D(n5647), .Z(
        n5622) );
  HS65_LS_AOI222X2 U13391 ( .A(n484), .B(n464), .C(n457), .D(n5646), .E(n479), 
        .F(n454), .Z(n5623) );
  HS65_LS_NAND4ABX3 U13392 ( .A(n7213), .B(n7214), .C(n7215), .D(n7216), .Z(
        n2818) );
  HS65_LS_CB4I6X4 U13393 ( .A(n301), .B(n300), .C(n281), .D(n7008), .Z(n7213)
         );
  HS65_LS_CBI4I1X3 U13394 ( .A(n6207), .B(n7157), .C(n7237), .D(n7239), .Z(
        n7214) );
  HS65_LS_AOI222X2 U13395 ( .A(n307), .B(n287), .C(n280), .D(n7238), .E(n302), 
        .F(n277), .Z(n7215) );
  HS65_LS_NAND4ABX3 U13396 ( .A(n7297), .B(n7298), .C(n7299), .D(n7300), .Z(
        n2776) );
  HS65_LS_OAI212X3 U13397 ( .A(n6081), .B(n6315), .C(n6312), .D(n6153), .E(
        n7355), .Z(n7298) );
  HS65_LS_NAND4ABX3 U13398 ( .A(n6654), .B(n6720), .C(n7357), .D(n7358), .Z(
        n7297) );
  HS65_LS_AOI212X2 U13399 ( .A(n551), .B(n563), .C(n571), .D(n547), .E(n7301), 
        .Z(n7300) );
  HS65_LS_NAND4ABX3 U13400 ( .A(n4732), .B(n4733), .C(n4734), .D(n4735), .Z(
        n2806) );
  HS65_LS_NAND4ABX3 U13401 ( .A(n4767), .B(n4768), .C(n4769), .D(n4770), .Z(
        n4732) );
  HS65_LS_OAI212X3 U13402 ( .A(n4759), .B(n4760), .C(n4464), .D(n4761), .E(
        n4762), .Z(n4733) );
  HS65_LS_AOI212X2 U13403 ( .A(n247), .B(n265), .C(n261), .D(n242), .E(n4736), 
        .Z(n4735) );
  HS65_LS_NAND4ABX3 U13404 ( .A(n4527), .B(n4528), .C(n4529), .D(n4530), .Z(
        n3543) );
  HS65_LS_CBI4I6X2 U13405 ( .A(n689), .B(n4531), .C(n695), .D(n4532), .Z(n4530) );
  HS65_LS_CBI4I1X3 U13406 ( .A(n4543), .B(n4544), .C(n4545), .D(n4546), .Z(
        n4527) );
  HS65_LS_AOI212X2 U13407 ( .A(n710), .B(n682), .C(n706), .D(n690), .E(n4536), 
        .Z(n4529) );
  HS65_LS_NAND4ABX3 U13408 ( .A(n6120), .B(n6121), .C(n6122), .D(n6123), .Z(
        n3218) );
  HS65_LS_CBI4I6X2 U13409 ( .A(n507), .B(n6124), .C(n513), .D(n6125), .Z(n6123) );
  HS65_LS_CBI4I1X3 U13410 ( .A(n6136), .B(n6137), .C(n6138), .D(n6139), .Z(
        n6120) );
  HS65_LS_AOI212X2 U13411 ( .A(n528), .B(n500), .C(n524), .D(n508), .E(n6129), 
        .Z(n6122) );
  HS65_LS_NAND4ABX3 U13412 ( .A(n5705), .B(n5706), .C(n5707), .D(n5708), .Z(
        n2784) );
  HS65_LS_OAI212X3 U13413 ( .A(n4488), .B(n4722), .C(n4719), .D(n4560), .E(
        n5763), .Z(n5706) );
  HS65_LS_NAND4ABX3 U13414 ( .A(n5061), .B(n5127), .C(n5765), .D(n5766), .Z(
        n5705) );
  HS65_LS_AOI212X2 U13415 ( .A(n25), .B(n37), .C(n45), .D(n21), .E(n5709), .Z(
        n5708) );
  HS65_LS_NAND4ABX3 U13416 ( .A(n5888), .B(n5889), .C(n5890), .D(n5891), .Z(
        n2825) );
  HS65_LS_MX41X4 U13417 ( .D0(n482), .S0(n462), .D1(n472), .S1(n453), .D2(n454), .S2(n483), .D3(n463), .S3(n4794), .Z(n5889) );
  HS65_LS_MX41X4 U13418 ( .D0(n481), .S0(n4616), .D1(n466), .S1(n477), .D2(
        n461), .S2(n471), .D3(n478), .S3(n457), .Z(n5888) );
  HS65_LS_NOR4ABX2 U13419 ( .A(n5405), .B(n5386), .C(n5892), .D(n4787), .Z(
        n5891) );
  HS65_LS_NAND4ABX3 U13420 ( .A(n7480), .B(n7481), .C(n7482), .D(n7483), .Z(
        n2817) );
  HS65_LS_MX41X4 U13421 ( .D0(n305), .S0(n285), .D1(n295), .S1(n276), .D2(n277), .S2(n306), .D3(n286), .S3(n6387), .Z(n7481) );
  HS65_LS_MX41X4 U13422 ( .D0(n304), .S0(n6209), .D1(n289), .S1(n300), .D2(
        n284), .S2(n294), .D3(n301), .S3(n280), .Z(n7480) );
  HS65_LS_NOR4ABX2 U13423 ( .A(n6997), .B(n6978), .C(n7484), .D(n6380), .Z(
        n7483) );
  HS65_LS_NAND4ABX3 U13424 ( .A(n7714), .B(n7715), .C(n7716), .D(n7717), .Z(
        n2809) );
  HS65_LS_NOR4ABX2 U13425 ( .A(n7718), .B(n7719), .C(n7720), .D(n7721), .Z(
        n7717) );
  HS65_LS_MX41X4 U13426 ( .D0(n126), .S0(n96), .D1(n110), .S1(n122), .D2(n107), 
        .S2(n127), .D3(n99), .S3(n7748), .Z(n7715) );
  HS65_LS_MX41X4 U13427 ( .D0(n128), .S0(n7747), .D1(n104), .S1(n138), .D2(n98), .S2(n124), .D3(n135), .S3(n113), .Z(n7714) );
  HS65_LS_NAND4ABX3 U13428 ( .A(n2836), .B(n2837), .C(n2838), .D(n2839), .Z(
        n2728) );
  HS65_LS_OAI212X3 U13429 ( .A(n2847), .B(n2848), .C(n2849), .D(n2850), .E(
        n2851), .Z(n2837) );
  HS65_LS_NAND4ABX3 U13430 ( .A(n2857), .B(n2858), .C(n2859), .D(n2860), .Z(
        n2836) );
  HS65_LS_AOI212X2 U13431 ( .A(n417), .B(n441), .C(n411), .D(n434), .E(n2840), 
        .Z(n2839) );
  HS65_LS_IVX2 U13432 ( .A(n3189), .Z(n430) );
  HS65_LS_NAND4ABX3 U13433 ( .A(n4771), .B(n4772), .C(n4773), .D(n4774), .Z(
        n2830) );
  HS65_LS_NAND4ABX3 U13434 ( .A(n4806), .B(n4807), .C(n4808), .D(n4809), .Z(
        n4771) );
  HS65_LS_OAI212X3 U13435 ( .A(n4798), .B(n4799), .C(n4510), .D(n4800), .E(
        n4801), .Z(n4772) );
  HS65_LS_AOI212X2 U13436 ( .A(n466), .B(n484), .C(n480), .D(n461), .E(n4775), 
        .Z(n4774) );
  HS65_LS_NAND4ABX3 U13437 ( .A(n3966), .B(n3967), .C(n3968), .D(n3969), .Z(
        n2717) );
  HS65_LS_CBI4I1X3 U13438 ( .A(n433), .B(n2847), .C(n3007), .D(n3986), .Z(
        n3967) );
  HS65_LS_AOI212X2 U13439 ( .A(n440), .B(n412), .C(n410), .D(n2861), .E(n3984), 
        .Z(n3968) );
  HS65_LS_CBI4I1X3 U13440 ( .A(n3209), .B(n2849), .C(n3004), .D(n3867), .Z(
        n3966) );
  HS65_LS_NAND4ABX3 U13441 ( .A(n3360), .B(n3361), .C(n3362), .D(n3363), .Z(
        n2707) );
  HS65_LS_OAI212X3 U13442 ( .A(n3413), .B(n2850), .C(n3414), .D(n3415), .E(
        n3416), .Z(n3361) );
  HS65_LS_NAND4ABX3 U13443 ( .A(n3417), .B(n3418), .C(n3419), .D(n3420), .Z(
        n3360) );
  HS65_LS_AOI212X2 U13444 ( .A(n410), .B(n3364), .C(n431), .D(n414), .E(n3365), 
        .Z(n3363) );
  HS65_LS_NAND4ABX3 U13445 ( .A(n2912), .B(n2913), .C(n2914), .D(n2915), .Z(
        n2640) );
  HS65_LS_CBI4I1X3 U13446 ( .A(n2923), .B(n2924), .C(n2925), .D(n2926), .Z(
        n2913) );
  HS65_LS_CBI4I1X3 U13447 ( .A(n2927), .B(n2928), .C(n2929), .D(n2930), .Z(
        n2912) );
  HS65_LS_AOI212X2 U13448 ( .A(n150), .B(n180), .C(n156), .D(n176), .E(n2921), 
        .Z(n2914) );
  HS65_LS_NAND4ABX3 U13449 ( .A(n2992), .B(n2993), .C(n2994), .D(n2995), .Z(
        n2696) );
  HS65_LS_CBI4I1X3 U13450 ( .A(n3007), .B(n2848), .C(n3008), .D(n3009), .Z(
        n2992) );
  HS65_LS_CBI4I1X3 U13451 ( .A(n3003), .B(n3004), .C(n3005), .D(n3006), .Z(
        n2993) );
  HS65_LS_AOI212X2 U13452 ( .A(n421), .B(n432), .C(n416), .D(n445), .E(n3001), 
        .Z(n2994) );
  HS65_LS_IVX2 U13453 ( .A(n8019), .Z(n390) );
  HS65_LS_IVX2 U13454 ( .A(n8061), .Z(n349) );
  HS65_LS_NAND4ABX3 U13455 ( .A(n6364), .B(n6365), .C(n6366), .D(n6367), .Z(
        n2822) );
  HS65_LS_NAND4ABX3 U13456 ( .A(n6399), .B(n6400), .C(n6401), .D(n6402), .Z(
        n6364) );
  HS65_LS_OAI212X3 U13457 ( .A(n6391), .B(n6392), .C(n6103), .D(n6393), .E(
        n6394), .Z(n6365) );
  HS65_LS_AOI212X2 U13458 ( .A(n289), .B(n307), .C(n303), .D(n284), .E(n6368), 
        .Z(n6367) );
  HS65_LS_NAND4ABX3 U13459 ( .A(n6407), .B(n6408), .C(n6409), .D(n6410), .Z(
        n3216) );
  HS65_LS_NAND4ABX3 U13460 ( .A(n6469), .B(n6470), .C(n6471), .D(n6472), .Z(
        n6407) );
  HS65_LS_OAI212X3 U13461 ( .A(n6465), .B(n6229), .C(n6466), .D(n6467), .E(
        n6468), .Z(n6408) );
  HS65_LS_AOI212X2 U13462 ( .A(n502), .B(n6411), .C(n530), .D(n505), .E(n6412), 
        .Z(n6410) );
  HS65_LS_NAND2X2 U13463 ( .A(n1469), .B(n1478), .Z(n1128) );
  HS65_LS_NAND2X2 U13464 ( .A(n2221), .B(n2230), .Z(n1880) );
  HS65_LS_NAND4ABX3 U13465 ( .A(n7421), .B(n7422), .C(n7423), .D(n7424), .Z(
        n2793) );
  HS65_LS_MX41X4 U13466 ( .D0(n84), .S0(n64), .D1(n74), .S1(n55), .D2(n56), 
        .S2(n85), .D3(n65), .S3(n6348), .Z(n7422) );
  HS65_LS_MX41X4 U13467 ( .D0(n83), .S0(n6184), .D1(n68), .S1(n79), .D2(n63), 
        .S2(n73), .D3(n80), .S3(n59), .Z(n7421) );
  HS65_LS_NOR4ABX2 U13468 ( .A(n6882), .B(n6863), .C(n7425), .D(n6341), .Z(
        n7424) );
  HS65_LS_NAND2X2 U13469 ( .A(n2597), .B(n2606), .Z(n2256) );
  HS65_LS_NAND2X2 U13470 ( .A(n1845), .B(n1854), .Z(n1504) );
  HS65_LS_NAND4ABX3 U13471 ( .A(n5829), .B(n5830), .C(n5831), .D(n5832), .Z(
        n2801) );
  HS65_LS_MX41X4 U13472 ( .D0(n263), .S0(n243), .D1(n253), .S1(n234), .D2(n235), .S2(n264), .D3(n244), .S3(n4755), .Z(n5830) );
  HS65_LS_MX41X4 U13473 ( .D0(n262), .S0(n4591), .D1(n247), .S1(n258), .D2(
        n242), .S2(n252), .D3(n259), .S3(n238), .Z(n5829) );
  HS65_LS_NOR4ABX2 U13474 ( .A(n5290), .B(n5271), .C(n5833), .D(n4748), .Z(
        n5832) );
  HS65_LS_NAND4ABX3 U13475 ( .A(n4814), .B(n4815), .C(n4816), .D(n4817), .Z(
        n3224) );
  HS65_LS_NAND4ABX3 U13476 ( .A(n4876), .B(n4877), .C(n4878), .D(n4879), .Z(
        n4814) );
  HS65_LS_OAI212X3 U13477 ( .A(n4872), .B(n4636), .C(n4873), .D(n4874), .E(
        n4875), .Z(n4815) );
  HS65_LS_AOI212X2 U13478 ( .A(n684), .B(n4818), .C(n712), .D(n687), .E(n4819), 
        .Z(n4817) );
  HS65_LS_NAND4ABX3 U13479 ( .A(n3916), .B(n3917), .C(n3918), .D(n3919), .Z(
        n2669) );
  HS65_LS_CBI4I1X3 U13480 ( .A(n3058), .B(n3262), .C(n2924), .D(n3634), .Z(
        n3916) );
  HS65_LS_CBI4I6X2 U13481 ( .A(n174), .B(n3608), .C(n159), .D(n3920), .Z(n3919) );
  HS65_LS_AOI212X2 U13482 ( .A(n172), .B(n157), .C(n158), .D(n3921), .E(n3922), 
        .Z(n3918) );
  HS65_LS_NAND4ABX3 U13483 ( .A(n8169), .B(n8170), .C(n8171), .D(n8172), .Z(
        n2814) );
  HS65_LS_NAND4ABX3 U13484 ( .A(n8197), .B(n8198), .C(n8199), .D(n8200), .Z(
        n8169) );
  HS65_LS_OAI212X3 U13485 ( .A(n7668), .B(n8192), .C(n7880), .D(n7917), .E(
        n8193), .Z(n8170) );
  HS65_LS_AOI212X2 U13486 ( .A(n104), .B(n125), .C(n137), .D(n98), .E(n8173), 
        .Z(n8172) );
  HS65_LS_NAND4ABX3 U13487 ( .A(n7652), .B(n7653), .C(n7654), .D(n7655), .Z(
        n2810) );
  HS65_LS_CBI4I1X3 U13488 ( .A(n7669), .B(n7666), .C(n7670), .D(n7671), .Z(
        n7653) );
  HS65_LS_CBI4I1X3 U13489 ( .A(n7672), .B(n7673), .C(n7674), .D(n7675), .Z(
        n7652) );
  HS65_LS_AOI222X2 U13490 ( .A(n125), .B(n97), .C(n113), .D(n7665), .E(n136), 
        .F(n107), .Z(n7654) );
  HS65_LS_NAND4ABX3 U13491 ( .A(n3230), .B(n3231), .C(n3232), .D(n3233), .Z(
        n2653) );
  HS65_LS_NAND4ABX3 U13492 ( .A(n3293), .B(n3294), .C(n3295), .D(n3296), .Z(
        n3230) );
  HS65_LS_OAI212X3 U13493 ( .A(n3289), .B(n3042), .C(n146), .D(n3290), .E(
        n3291), .Z(n3231) );
  HS65_LS_AOI212X2 U13494 ( .A(n158), .B(n3234), .C(n182), .D(n153), .E(n3235), 
        .Z(n3233) );
  HS65_LS_NAND4ABX3 U13495 ( .A(n7166), .B(n7167), .C(n7168), .D(n7169), .Z(
        n3017) );
  HS65_LS_CB4I6X4 U13496 ( .A(n515), .B(n514), .C(n501), .D(n6777), .Z(n7166)
         );
  HS65_LS_CBI4I1X3 U13497 ( .A(n6138), .B(n7181), .C(n7183), .D(n7185), .Z(
        n7167) );
  HS65_LS_AOI222X2 U13498 ( .A(n517), .B(n498), .C(n502), .D(n7184), .E(n511), 
        .F(n506), .Z(n7168) );
  HS65_LS_NAND4ABX3 U13499 ( .A(n5574), .B(n5575), .C(n5576), .D(n5577), .Z(
        n3221) );
  HS65_LS_CB4I6X4 U13500 ( .A(n697), .B(n696), .C(n683), .D(n5185), .Z(n5574)
         );
  HS65_LS_CBI4I1X3 U13501 ( .A(n4545), .B(n5589), .C(n5591), .D(n5593), .Z(
        n5575) );
  HS65_LS_AOI222X2 U13502 ( .A(n699), .B(n680), .C(n684), .D(n5592), .E(n693), 
        .F(n688), .Z(n5576) );
  HS65_LS_NAND4ABX3 U13503 ( .A(n4030), .B(n4031), .C(n4032), .D(n4033), .Z(
        n2722) );
  HS65_LS_CB4I6X4 U13504 ( .A(n436), .B(n435), .C(n412), .D(n3860), .Z(n4030)
         );
  HS65_LS_AOI222X2 U13505 ( .A(n422), .B(n442), .C(n410), .D(n4052), .E(n415), 
        .F(n438), .Z(n4032) );
  HS65_LS_CBI4I1X3 U13506 ( .A(n3008), .B(n3214), .C(n3895), .D(n4053), .Z(
        n4031) );
  HS65_LS_NAND4ABX3 U13507 ( .A(n3134), .B(n3135), .C(n3136), .D(n3137), .Z(
        n2647) );
  HS65_LS_NAND4ABX3 U13508 ( .A(n3169), .B(n3170), .C(n3171), .D(n3172), .Z(
        n3134) );
  HS65_LS_OAI212X3 U13509 ( .A(n3161), .B(n3162), .C(n3163), .D(n2893), .E(
        n3164), .Z(n3135) );
  HS65_LS_AOI212X2 U13510 ( .A(n648), .B(n666), .C(n643), .D(n661), .E(n3138), 
        .Z(n3137) );
  HS65_LS_NAND4ABX3 U13511 ( .A(n3928), .B(n3929), .C(n3930), .D(n3931), .Z(
        n2681) );
  HS65_LS_CB4I6X4 U13512 ( .A(n214), .B(n213), .C(n202), .D(n3502), .Z(n3928)
         );
  HS65_LS_CBI4I1X3 U13513 ( .A(n2879), .B(n2971), .C(n3538), .D(n3944), .Z(
        n3929) );
  HS65_LS_AOI222X2 U13514 ( .A(n194), .B(n215), .C(n203), .D(n3943), .E(n199), 
        .F(n210), .Z(n3930) );
  HS65_LS_NAND4ABX3 U13515 ( .A(n9063), .B(n9064), .C(n9065), .D(n9066), .Z(
        n2811) );
  HS65_LS_CBI4I1X3 U13516 ( .A(n120), .B(n7725), .C(n7735), .D(n9120), .Z(
        n9064) );
  HS65_LS_AOI212X2 U13517 ( .A(n112), .B(n126), .C(n113), .D(n7891), .E(n9118), 
        .Z(n9065) );
  HS65_LS_CBI4I1X3 U13518 ( .A(n7672), .B(n7881), .C(n8472), .D(n8801), .Z(
        n9063) );
  HS65_LS_NAND4ABX3 U13519 ( .A(n5550), .B(n5551), .C(n5552), .D(n5553), .Z(
        n2827) );
  HS65_LS_AOI212X2 U13520 ( .A(n458), .B(n482), .C(n457), .D(n4523), .E(n5569), 
        .Z(n5552) );
  HS65_LS_CBI4I1X3 U13521 ( .A(n4805), .B(n4512), .C(n4989), .D(n5413), .Z(
        n5550) );
  HS65_LS_CBI4I1X3 U13522 ( .A(n476), .B(n4509), .C(n4613), .D(n5570), .Z(
        n5551) );
  HS65_LS_NAND4ABX3 U13523 ( .A(n7142), .B(n7143), .C(n7144), .D(n7145), .Z(
        n2819) );
  HS65_LS_AOI212X2 U13524 ( .A(n281), .B(n305), .C(n280), .D(n6116), .E(n7161), 
        .Z(n7144) );
  HS65_LS_CBI4I1X3 U13525 ( .A(n6398), .B(n6105), .C(n6582), .D(n7005), .Z(
        n7142) );
  HS65_LS_CBI4I1X3 U13526 ( .A(n299), .B(n6102), .C(n6206), .D(n7162), .Z(
        n7143) );
  HS65_LS_IVX2 U13527 ( .A(n7857), .Z(n365) );
  HS65_LS_NAND4ABX3 U13528 ( .A(n6325), .B(n6326), .C(n6327), .D(n6328), .Z(
        n2798) );
  HS65_LS_NAND4ABX3 U13529 ( .A(n6360), .B(n6361), .C(n6362), .D(n6363), .Z(
        n6325) );
  HS65_LS_OAI212X3 U13530 ( .A(n6352), .B(n6353), .C(n6057), .D(n6354), .E(
        n6355), .Z(n6326) );
  HS65_LS_AOI212X2 U13531 ( .A(n68), .B(n86), .C(n82), .D(n63), .E(n6329), .Z(
        n6328) );
  HS65_LS_NAND4ABX3 U13532 ( .A(n8944), .B(n8945), .C(n8946), .D(n8947), .Z(
        n2762) );
  HS65_LS_CBI4I1X3 U13533 ( .A(n7863), .B(n7871), .C(n7761), .D(n9004), .Z(
        n8945) );
  HS65_LS_AOI222X2 U13534 ( .A(n372), .B(n397), .C(n376), .D(n9003), .E(n403), 
        .F(n378), .Z(n8946) );
  HS65_LS_CBI4I1X3 U13535 ( .A(n7869), .B(n8663), .C(n8004), .D(n8284), .Z(
        n8944) );
  HS65_LS_NAND2X2 U13536 ( .A(n4339), .B(n4340), .Z(n2848) );
  HS65_LS_NAND4ABX3 U13537 ( .A(n3945), .B(n3946), .C(n3947), .D(n3948), .Z(
        n2667) );
  HS65_LS_AOI212X2 U13538 ( .A(n664), .B(n635), .C(n633), .D(n2906), .E(n3963), 
        .Z(n3947) );
  HS65_LS_CBI4I1X3 U13539 ( .A(n657), .B(n2892), .C(n2989), .D(n3965), .Z(
        n3946) );
  HS65_LS_CBI4I1X3 U13540 ( .A(n3168), .B(n2894), .C(n2986), .D(n3750), .Z(
        n3945) );
  HS65_LS_IVX2 U13541 ( .A(n2946), .Z(n227) );
  HS65_LS_IVX2 U13542 ( .A(n3148), .Z(n654) );
  HS65_LS_NOR4ABX2 U13543 ( .A(n3970), .B(n3971), .C(n3972), .D(n3973), .Z(
        n3969) );
  HS65_LS_OAI212X3 U13544 ( .A(n3415), .B(n3895), .C(n3189), .D(n2850), .E(
        n2844), .Z(n3972) );
  HS65_LS_NAND4ABX3 U13545 ( .A(n4547), .B(n4548), .C(n4549), .D(n4550), .Z(
        n2782) );
  HS65_LS_NAND4ABX3 U13546 ( .A(n4583), .B(n4584), .C(n4585), .D(n4586), .Z(
        n4547) );
  HS65_LS_OAI212X3 U13547 ( .A(n4575), .B(n4576), .C(n4488), .D(n4577), .E(
        n4578), .Z(n4548) );
  HS65_LS_AOI212X2 U13548 ( .A(n10), .B(n35), .C(n31), .D(n14), .E(n4551), .Z(
        n4550) );
  HS65_LS_NAND4ABX3 U13549 ( .A(n6140), .B(n6141), .C(n6142), .D(n6143), .Z(
        n2774) );
  HS65_LS_NAND4ABX3 U13550 ( .A(n6176), .B(n6177), .C(n6178), .D(n6179), .Z(
        n6140) );
  HS65_LS_OAI212X3 U13551 ( .A(n6168), .B(n6169), .C(n6081), .D(n6170), .E(
        n6171), .Z(n6141) );
  HS65_LS_AOI212X2 U13552 ( .A(n536), .B(n561), .C(n557), .D(n540), .E(n6144), 
        .Z(n6143) );
  HS65_LS_NAND2X2 U13553 ( .A(n9053), .B(n9030), .Z(n7817) );
  HS65_LS_NAND2X2 U13554 ( .A(n9111), .B(n9088), .Z(n7880) );
  HS65_LS_NAND4ABX3 U13555 ( .A(n5480), .B(n5481), .C(n5482), .D(n5483), .Z(
        n2779) );
  HS65_LS_CBI4I1X3 U13556 ( .A(n4582), .B(n4719), .C(n4720), .D(n5059), .Z(
        n5480) );
  HS65_LS_AOI212X2 U13557 ( .A(n18), .B(n38), .C(n20), .D(n5489), .E(n5490), 
        .Z(n5482) );
  HS65_LS_CBI4I1X3 U13558 ( .A(n30), .B(n4722), .C(n4487), .D(n5491), .Z(n5481) );
  HS65_LS_NAND4ABX3 U13559 ( .A(n7072), .B(n7073), .C(n7074), .D(n7075), .Z(
        n2771) );
  HS65_LS_CBI4I1X3 U13560 ( .A(n6175), .B(n6312), .C(n6313), .D(n6652), .Z(
        n7072) );
  HS65_LS_AOI212X2 U13561 ( .A(n544), .B(n564), .C(n546), .D(n7081), .E(n7082), 
        .Z(n7074) );
  HS65_LS_CBI4I1X3 U13562 ( .A(n556), .B(n6315), .C(n6080), .D(n7083), .Z(
        n7073) );
  HS65_LS_NAND4ABX3 U13563 ( .A(n8384), .B(n8385), .C(n8386), .D(n8387), .Z(
        n2789) );
  HS65_LS_NAND4ABX3 U13564 ( .A(n8432), .B(n8433), .C(n8434), .D(n8435), .Z(
        n8384) );
  HS65_LS_OAI212X3 U13565 ( .A(n8430), .B(n7632), .C(n590), .D(n7639), .E(
        n8431), .Z(n8385) );
  HS65_LS_AOI212X2 U13566 ( .A(n600), .B(n8388), .C(n597), .D(n609), .E(n8389), 
        .Z(n8387) );
  HS65_LS_NAND4ABX3 U13567 ( .A(n7101), .B(n7102), .C(n7103), .D(n7104), .Z(
        n2770) );
  HS65_LS_CB4I6X4 U13568 ( .A(n559), .B(n558), .C(n544), .D(n6656), .Z(n7101)
         );
  HS65_LS_CBI4I1X3 U13569 ( .A(n6082), .B(n7116), .C(n7118), .D(n7120), .Z(
        n7102) );
  HS65_LS_AOI222X2 U13570 ( .A(n541), .B(n561), .C(n546), .D(n7119), .E(n550), 
        .F(n555), .Z(n7103) );
  HS65_LS_NAND4ABX3 U13571 ( .A(n5509), .B(n5510), .C(n5511), .D(n5512), .Z(
        n2778) );
  HS65_LS_CB4I6X4 U13572 ( .A(n33), .B(n32), .C(n18), .D(n5063), .Z(n5509) );
  HS65_LS_CBI4I1X3 U13573 ( .A(n4489), .B(n5524), .C(n5526), .D(n5528), .Z(
        n5510) );
  HS65_LS_AOI222X2 U13574 ( .A(n15), .B(n35), .C(n20), .D(n5527), .E(n24), .F(
        n29), .Z(n5511) );
  HS65_LS_IVX2 U13575 ( .A(n1529), .Z(n833) );
  HS65_LS_IVX2 U13576 ( .A(n2281), .Z(n915) );
  HS65_LS_IVX2 U13577 ( .A(n1153), .Z(n874) );
  HS65_LS_IVX2 U13578 ( .A(n1905), .Z(n792) );
  HS65_LS_OAI212X3 U13579 ( .A(n4188), .B(n3470), .C(n3484), .D(n3454), .E(
        n4189), .Z(n4187) );
  HS65_LS_OAI21X2 U13580 ( .A(n200), .B(n195), .C(n221), .Z(n4189) );
  HS65_LS_NOR3X1 U13581 ( .A(n215), .B(n225), .C(n227), .Z(n4188) );
  HS65_LS_IVX2 U13582 ( .A(n1879), .Z(n778) );
  HS65_LS_IVX2 U13583 ( .A(n1503), .Z(n819) );
  HS65_LS_IVX2 U13584 ( .A(n2255), .Z(n901) );
  HS65_LS_IVX2 U13585 ( .A(n1127), .Z(n860) );
  HS65_LS_NAND4ABX3 U13586 ( .A(n7624), .B(n7625), .C(n7626), .D(n7627), .Z(
        n2786) );
  HS65_LS_CBI4I1X3 U13587 ( .A(n7641), .B(n7638), .C(n7642), .D(n7643), .Z(
        n7625) );
  HS65_LS_CBI4I1X3 U13588 ( .A(n7644), .B(n7645), .C(n7646), .D(n7647), .Z(
        n7624) );
  HS65_LS_AOI222X2 U13589 ( .A(n612), .B(n584), .C(n600), .D(n7637), .E(n623), 
        .F(n594), .Z(n7626) );
  HS65_LS_IVX2 U13590 ( .A(n8436), .Z(n624) );
  HS65_LS_IVX2 U13591 ( .A(n8447), .Z(n137) );
  HS65_LS_NAND2X2 U13592 ( .A(n8935), .B(n8928), .Z(n7964) );
  HS65_LS_IVX2 U13593 ( .A(n3625), .Z(n160) );
  HS65_LS_IVX2 U13594 ( .A(n3454), .Z(n203) );
  HS65_LS_IVX2 U13595 ( .A(n2984), .Z(n633) );
  HS65_LS_IVX2 U13596 ( .A(n3002), .Z(n410) );
  HS65_LS_IVX2 U13597 ( .A(n2847), .Z(n443) );
  HS65_LS_NAND2X2 U13598 ( .A(n4280), .B(n4281), .Z(n2893) );
  HS65_LS_IVX2 U13599 ( .A(n5645), .Z(n461) );
  HS65_LS_IVX2 U13600 ( .A(n5618), .Z(n242) );
  HS65_LS_IVX2 U13601 ( .A(n7237), .Z(n284) );
  HS65_LS_IVX2 U13602 ( .A(n7210), .Z(n63) );
  HS65_LS_IVX2 U13603 ( .A(n5591), .Z(n679) );
  HS65_LS_IVX2 U13604 ( .A(n7183), .Z(n497) );
  HS65_LS_IVX2 U13605 ( .A(n2892), .Z(n667) );
  HS65_LS_NAND4ABX3 U13606 ( .A(n5594), .B(n5595), .C(n5596), .D(n5597), .Z(
        n2802) );
  HS65_LS_CB4I6X4 U13607 ( .A(n259), .B(n258), .C(n239), .D(n5301), .Z(n5594)
         );
  HS65_LS_CBI4I1X3 U13608 ( .A(n4602), .B(n5544), .C(n5618), .D(n5620), .Z(
        n5595) );
  HS65_LS_AOI222X2 U13609 ( .A(n265), .B(n245), .C(n238), .D(n5619), .E(n260), 
        .F(n235), .Z(n5596) );
  HS65_LS_IVX2 U13610 ( .A(n3102), .Z(n219) );
  HS65_LS_IVX2 U13611 ( .A(n6270), .Z(n557) );
  HS65_LS_IVX2 U13612 ( .A(n4677), .Z(n31) );
  HS65_LS_IVX2 U13613 ( .A(n4881), .Z(n695) );
  HS65_LS_IVX2 U13614 ( .A(n5009), .Z(n480) );
  HS65_LS_IVX2 U13615 ( .A(n6602), .Z(n303) );
  HS65_LS_IVX2 U13616 ( .A(n6488), .Z(n82) );
  HS65_LS_IVX2 U13617 ( .A(n6474), .Z(n513) );
  HS65_LS_IVX2 U13618 ( .A(n4895), .Z(n261) );
  HS65_LS_IVX2 U13619 ( .A(n4509), .Z(n487) );
  HS65_LS_IVX2 U13620 ( .A(n4463), .Z(n268) );
  HS65_LS_IVX2 U13621 ( .A(n6102), .Z(n310) );
  HS65_LS_IVX2 U13622 ( .A(n6056), .Z(n89) );
  HS65_LS_IVX2 U13623 ( .A(n4862), .Z(n704) );
  HS65_LS_IVX2 U13624 ( .A(n6455), .Z(n522) );
  HS65_LS_NAND4ABX3 U13625 ( .A(n4498), .B(n4499), .C(n4500), .D(n4501), .Z(
        n2832) );
  HS65_LS_NAND4ABX3 U13626 ( .A(n4519), .B(n4520), .C(n4521), .D(n4522), .Z(
        n4498) );
  HS65_LS_OAI212X3 U13627 ( .A(n4509), .B(n4510), .C(n4511), .D(n4512), .E(
        n4513), .Z(n4499) );
  HS65_LS_AOI212X2 U13628 ( .A(n455), .B(n483), .C(n459), .D(n475), .E(n4502), 
        .Z(n4501) );
  HS65_LS_NAND4ABX3 U13629 ( .A(n6091), .B(n6092), .C(n6093), .D(n6094), .Z(
        n2824) );
  HS65_LS_NAND4ABX3 U13630 ( .A(n6112), .B(n6113), .C(n6114), .D(n6115), .Z(
        n6091) );
  HS65_LS_OAI212X3 U13631 ( .A(n6102), .B(n6103), .C(n6104), .D(n6105), .E(
        n6106), .Z(n6092) );
  HS65_LS_AOI212X2 U13632 ( .A(n278), .B(n306), .C(n282), .D(n298), .E(n6095), 
        .Z(n6094) );
  HS65_LS_IVX2 U13633 ( .A(n3290), .Z(n180) );
  HS65_LS_IVX2 U13634 ( .A(n4874), .Z(n710) );
  HS65_LS_IVX2 U13635 ( .A(n5002), .Z(n474) );
  HS65_LS_IVX2 U13636 ( .A(n6595), .Z(n297) );
  HS65_LS_IVX2 U13637 ( .A(n6481), .Z(n76) );
  HS65_LS_IVX2 U13638 ( .A(n6467), .Z(n528) );
  HS65_LS_IVX2 U13639 ( .A(n4888), .Z(n255) );
  HS65_LS_IVX2 U13640 ( .A(n5026), .Z(n20) );
  HS65_LS_IVX2 U13641 ( .A(n6619), .Z(n546) );
  HS65_LS_IVX2 U13642 ( .A(n4620), .Z(n457) );
  HS65_LS_IVX2 U13643 ( .A(n4595), .Z(n238) );
  HS65_LS_IVX2 U13644 ( .A(n6213), .Z(n280) );
  HS65_LS_IVX2 U13645 ( .A(n6188), .Z(n59) );
  HS65_LS_IVX2 U13646 ( .A(n5148), .Z(n684) );
  HS65_LS_IVX2 U13647 ( .A(n6740), .Z(n502) );
  HS65_LS_IVX2 U13648 ( .A(n2336), .Z(n894) );
  HS65_LS_IVX2 U13649 ( .A(n1584), .Z(n812) );
  HS65_LS_IVX2 U13650 ( .A(n1201), .Z(n858) );
  HS65_LS_IVX2 U13651 ( .A(n1953), .Z(n776) );
  HS65_LS_IVX2 U13652 ( .A(n1577), .Z(n817) );
  HS65_LS_IVX2 U13653 ( .A(n2329), .Z(n899) );
  HS65_LS_IVX2 U13654 ( .A(n1208), .Z(n853) );
  HS65_LS_IVX2 U13655 ( .A(n1960), .Z(n771) );
  HS65_LS_IVX2 U13656 ( .A(n6262), .Z(n572) );
  HS65_LS_IVX2 U13657 ( .A(n4669), .Z(n46) );
  HS65_LS_IVX2 U13658 ( .A(n3168), .Z(n660) );
  HS65_LS_IVX2 U13659 ( .A(n5526), .Z(n14) );
  HS65_LS_IVX2 U13660 ( .A(n7118), .Z(n540) );
  HS65_LS_IVX2 U13661 ( .A(n3599), .Z(n158) );
  HS65_LS_IVX2 U13662 ( .A(n7832), .Z(n600) );
  HS65_LS_IVX2 U13663 ( .A(n7931), .Z(n113) );
  HS65_LS_OAI212X3 U13664 ( .A(n610), .B(n7686), .C(n8436), .D(n8159), .E(
        n9043), .Z(n9041) );
  HS65_LS_IVX2 U13665 ( .A(n8750), .Z(n610) );
  HS65_LS_CBI4I6X2 U13666 ( .A(n623), .B(n615), .C(n601), .D(n8748), .Z(n9043)
         );
  HS65_LS_OAI212X3 U13667 ( .A(n123), .B(n7724), .C(n8447), .D(n8191), .E(
        n9101), .Z(n9099) );
  HS65_LS_IVX2 U13668 ( .A(n8838), .Z(n123) );
  HS65_LS_CBI4I6X2 U13669 ( .A(n136), .B(n128), .C(n114), .D(n8836), .Z(n9101)
         );
  HS65_LS_IVX2 U13670 ( .A(n7672), .Z(n135) );
  HS65_LS_IVX2 U13671 ( .A(n7644), .Z(n622) );
  HS65_LS_IVX2 U13672 ( .A(n8412), .Z(n593) );
  HS65_LS_IVX2 U13673 ( .A(n8472), .Z(n106) );
  HS65_LS_NAND4ABX3 U13674 ( .A(n8626), .B(n8627), .C(n8628), .D(n8629), .Z(
        n3015) );
  HS65_LS_OAI212X3 U13675 ( .A(n7964), .B(n7779), .C(n8361), .D(n7955), .E(
        n8640), .Z(n8627) );
  HS65_LS_NAND4ABX3 U13676 ( .A(n8642), .B(n8538), .C(n8579), .D(n8643), .Z(
        n8626) );
  HS65_LS_AOI212X2 U13677 ( .A(n332), .B(n353), .C(n327), .D(n348), .E(n8630), 
        .Z(n8629) );
  HS65_LS_IVX2 U13678 ( .A(n3264), .Z(n174) );
  HS65_LS_IVX2 U13679 ( .A(n7952), .Z(n344) );
  HS65_LS_IVX2 U13680 ( .A(n8220), .Z(n376) );
  HS65_LS_NAND2X2 U13681 ( .A(n4147), .B(n4162), .Z(n2928) );
  HS65_LS_IVX2 U13682 ( .A(n2966), .Z(n214) );
  HS65_LS_IVX2 U13683 ( .A(n3209), .Z(n436) );
  HS65_LS_IVX2 U13684 ( .A(n3895), .Z(n419) );
  HS65_LS_IVX2 U13685 ( .A(n3470), .Z(n189) );
  HS65_LS_IVX2 U13686 ( .A(n4103), .Z(n165) );
  HS65_LS_IVX2 U13687 ( .A(n7639), .Z(n608) );
  HS65_LS_IVX2 U13688 ( .A(n7667), .Z(n121) );
  HS65_LS_IVX2 U13689 ( .A(n3353), .Z(n656) );
  HS65_LS_OAI212X3 U13690 ( .A(n34), .B(n4680), .C(n4721), .D(n4677), .E(n5525), .Z(n5521) );
  HS65_LS_IVX2 U13691 ( .A(n5125), .Z(n34) );
  HS65_LS_CBI4I6X2 U13692 ( .A(n29), .B(n36), .C(n21), .D(n5118), .Z(n5525) );
  HS65_LS_OAI212X3 U13693 ( .A(n560), .B(n6273), .C(n6314), .D(n6270), .E(
        n7117), .Z(n7113) );
  HS65_LS_IVX2 U13694 ( .A(n6718), .Z(n560) );
  HS65_LS_CBI4I6X2 U13695 ( .A(n555), .B(n562), .C(n547), .D(n6711), .Z(n7117)
         );
  HS65_LS_NAND4ABX3 U13696 ( .A(n8137), .B(n8138), .C(n8139), .D(n8140), .Z(
        n2790) );
  HS65_LS_NAND4ABX3 U13697 ( .A(n8165), .B(n8166), .C(n8167), .D(n8168), .Z(
        n8137) );
  HS65_LS_OAI212X3 U13698 ( .A(n7640), .B(n8160), .C(n7817), .D(n7818), .E(
        n8161), .Z(n8138) );
  HS65_LS_AOI212X2 U13699 ( .A(n591), .B(n612), .C(n624), .D(n585), .E(n8141), 
        .Z(n8140) );
  HS65_LS_OAI212X3 U13700 ( .A(n8569), .B(n8070), .C(n7961), .D(n7964), .E(
        n8570), .Z(n8559) );
  HS65_LS_NOR2X2 U13701 ( .A(n337), .B(n8513), .Z(n8569) );
  HS65_LS_OAI212X3 U13702 ( .A(n3623), .B(n3280), .C(n2925), .D(n2928), .E(
        n3624), .Z(n3613) );
  HS65_LS_NOR2X2 U13703 ( .A(n152), .B(n3552), .Z(n3623) );
  HS65_LS_OAI212X3 U13704 ( .A(n8316), .B(n7760), .C(n7859), .D(n8030), .E(
        n8986), .Z(n8984) );
  HS65_LS_CB4I1X4 U13705 ( .A(n8671), .B(n8009), .C(n8267), .D(n8317), .Z(
        n8986) );
  HS65_LS_IVX2 U13706 ( .A(n6186), .Z(n81) );
  HS65_LS_IVX2 U13707 ( .A(n4618), .Z(n479) );
  HS65_LS_IVX2 U13708 ( .A(n6211), .Z(n302) );
  HS65_LS_IVX2 U13709 ( .A(n4593), .Z(n260) );
  HS65_LS_IVX2 U13710 ( .A(n4534), .Z(n693) );
  HS65_LS_IVX2 U13711 ( .A(n6127), .Z(n511) );
  HS65_LS_NAND4ABX3 U13712 ( .A(n3298), .B(n3299), .C(n3300), .D(n3301), .Z(
        n2745) );
  HS65_LS_OAI212X3 U13713 ( .A(n3351), .B(n2895), .C(n3352), .D(n3353), .E(
        n3354), .Z(n3299) );
  HS65_LS_NAND4ABX3 U13714 ( .A(n3355), .B(n3356), .C(n3357), .D(n3358), .Z(
        n3298) );
  HS65_LS_AOI212X2 U13715 ( .A(n633), .B(n3302), .C(n655), .D(n637), .E(n3303), 
        .Z(n3301) );
  HS65_LS_IVX2 U13716 ( .A(n7869), .Z(n401) );
  HS65_LS_IVX2 U13717 ( .A(n4805), .Z(n478) );
  HS65_LS_IVX2 U13718 ( .A(n6398), .Z(n301) );
  HS65_LS_IVX2 U13719 ( .A(n6359), .Z(n80) );
  HS65_LS_IVX2 U13720 ( .A(n4766), .Z(n259) );
  HS65_LS_IVX2 U13721 ( .A(n4659), .Z(n697) );
  HS65_LS_IVX2 U13722 ( .A(n6252), .Z(n515) );
  HS65_LS_IVX2 U13723 ( .A(n3063), .Z(n143) );
  HS65_LS_IVX2 U13724 ( .A(n3058), .Z(n168) );
  HS65_LS_IVX2 U13725 ( .A(n4582), .Z(n33) );
  HS65_LS_IVX2 U13726 ( .A(n6175), .Z(n559) );
  HS65_LS_NAND4ABX3 U13727 ( .A(n9005), .B(n9006), .C(n9007), .D(n9008), .Z(
        n2787) );
  HS65_LS_CBI4I1X3 U13728 ( .A(n607), .B(n7687), .C(n7697), .D(n9062), .Z(
        n9006) );
  HS65_LS_AOI212X2 U13729 ( .A(n599), .B(n613), .C(n600), .D(n7852), .E(n9060), 
        .Z(n9007) );
  HS65_LS_CBI4I1X3 U13730 ( .A(n7644), .B(n7842), .C(n8412), .D(n8713), .Z(
        n9005) );
  HS65_LS_NAND4ABX3 U13731 ( .A(n7121), .B(n7122), .C(n7123), .D(n7124), .Z(
        n2795) );
  HS65_LS_AOI212X2 U13732 ( .A(n60), .B(n84), .C(n59), .D(n6070), .E(n7140), 
        .Z(n7123) );
  HS65_LS_CBI4I1X3 U13733 ( .A(n6359), .B(n6059), .C(n6528), .D(n6890), .Z(
        n7121) );
  HS65_LS_CBI4I1X3 U13734 ( .A(n78), .B(n6056), .C(n6194), .D(n7141), .Z(n7122) );
  HS65_LS_NAND4ABX3 U13735 ( .A(n5529), .B(n5530), .C(n5531), .D(n5532), .Z(
        n2803) );
  HS65_LS_AOI212X2 U13736 ( .A(n239), .B(n263), .C(n238), .D(n4477), .E(n5548), 
        .Z(n5531) );
  HS65_LS_CBI4I1X3 U13737 ( .A(n4766), .B(n4466), .C(n4935), .D(n5298), .Z(
        n5529) );
  HS65_LS_CBI4I1X3 U13738 ( .A(n257), .B(n4463), .C(n4601), .D(n5549), .Z(
        n5530) );
  HS65_LS_IVX2 U13739 ( .A(n6087), .Z(n555) );
  HS65_LS_IVX2 U13740 ( .A(n4494), .Z(n29) );
  HS65_LS_NOR4ABX2 U13741 ( .A(n7948), .B(n7949), .C(n7950), .D(n7951), .Z(
        n7947) );
  HS65_LS_OAI212X3 U13742 ( .A(n7952), .B(n7953), .C(n7954), .D(n7955), .E(
        n7956), .Z(n7950) );
  HS65_LS_OAI212X3 U13743 ( .A(n3042), .B(n3043), .C(n3044), .D(n3045), .E(
        n3046), .Z(n3032) );
  HS65_LS_OAI21X2 U13744 ( .A(n160), .B(n159), .C(n174), .Z(n3046) );
  HS65_LS_OAI212X3 U13745 ( .A(n8094), .B(n8095), .C(n7998), .D(n8080), .E(
        n8096), .Z(n8083) );
  HS65_LS_OAI21X2 U13746 ( .A(n375), .B(n369), .C(n399), .Z(n8096) );
  HS65_LS_NOR2X2 U13747 ( .A(n378), .B(n380), .Z(n8094) );
  HS65_LS_IVX2 U13748 ( .A(n7991), .Z(n136) );
  HS65_LS_IVX2 U13749 ( .A(n7978), .Z(n623) );
  HS65_LS_IVX2 U13750 ( .A(n3726), .Z(n665) );
  HS65_LS_IVX2 U13751 ( .A(n3843), .Z(n441) );
  HS65_LS_IVX2 U13752 ( .A(n3484), .Z(n216) );
  HS65_LS_OAI212X3 U13753 ( .A(n3725), .B(n3726), .C(n2987), .D(n2893), .E(
        n3727), .Z(n3715) );
  HS65_LS_NOR2X2 U13754 ( .A(n644), .B(n3670), .Z(n3725) );
  HS65_LS_IVX2 U13755 ( .A(n5566), .Z(n481) );
  HS65_LS_IVX2 U13756 ( .A(n5545), .Z(n262) );
  HS65_LS_IVX2 U13757 ( .A(n5581), .Z(n700) );
  HS65_LS_IVX2 U13758 ( .A(n7158), .Z(n304) );
  HS65_LS_IVX2 U13759 ( .A(n7137), .Z(n83) );
  HS65_LS_IVX2 U13760 ( .A(n7173), .Z(n518) );
  HS65_LS_IVX2 U13761 ( .A(n8671), .Z(n403) );
  HS65_LS_OAI212X3 U13762 ( .A(n2437), .B(n2438), .C(n2284), .D(n2256), .E(
        n2439), .Z(n2427) );
  HS65_LS_NOR2X2 U13763 ( .A(n924), .B(n2398), .Z(n2437) );
  HS65_LS_OAI212X3 U13764 ( .A(n1685), .B(n1686), .C(n1532), .D(n1504), .E(
        n1687), .Z(n1675) );
  HS65_LS_NOR2X2 U13765 ( .A(n842), .B(n1646), .Z(n1685) );
  HS65_LS_OAI212X3 U13766 ( .A(n1309), .B(n1310), .C(n1156), .D(n1128), .E(
        n1311), .Z(n1299) );
  HS65_LS_NOR2X2 U13767 ( .A(n883), .B(n1270), .Z(n1309) );
  HS65_LS_OAI212X3 U13768 ( .A(n8265), .B(n8031), .C(n7859), .D(n7862), .E(
        n8266), .Z(n8255) );
  HS65_LS_NOR2X2 U13769 ( .A(n371), .B(n8208), .Z(n8265) );
  HS65_LS_IVX2 U13770 ( .A(n7084), .Z(n541) );
  HS65_LS_IVX2 U13771 ( .A(n5492), .Z(n15) );
  HS65_LS_IVX2 U13772 ( .A(n5516), .Z(n36) );
  HS65_LS_IVX2 U13773 ( .A(n7108), .Z(n562) );
  HS65_LS_OAI212X3 U13774 ( .A(n2061), .B(n2062), .C(n1908), .D(n1880), .E(
        n2063), .Z(n2051) );
  HS65_LS_NOR2X2 U13775 ( .A(n801), .B(n2022), .Z(n2061) );
  HS65_LS_IVX2 U13776 ( .A(n4002), .Z(n167) );
  HS65_LS_IVX2 U13777 ( .A(n1404), .Z(n854) );
  HS65_LS_IVX2 U13778 ( .A(n2156), .Z(n772) );
  HS65_LS_IVX2 U13779 ( .A(n1780), .Z(n813) );
  HS65_LS_IVX2 U13780 ( .A(n2532), .Z(n895) );
  HS65_LS_IVX2 U13781 ( .A(n1130), .Z(n889) );
  HS65_LS_IVX2 U13782 ( .A(n1882), .Z(n807) );
  HS65_LS_IVX2 U13783 ( .A(n1506), .Z(n848) );
  HS65_LS_IVX2 U13784 ( .A(n2258), .Z(n930) );
  HS65_LS_IVX2 U13785 ( .A(n6064), .Z(n66) );
  HS65_LS_IVX2 U13786 ( .A(n4517), .Z(n464) );
  HS65_LS_IVX2 U13787 ( .A(n6110), .Z(n287) );
  HS65_LS_IVX2 U13788 ( .A(n4471), .Z(n245) );
  HS65_LS_IVX2 U13789 ( .A(n5508), .Z(n680) );
  HS65_LS_IVX2 U13790 ( .A(n7100), .Z(n498) );
  HS65_LS_IVX2 U13791 ( .A(n8080), .Z(n394) );
  HS65_LS_IVX2 U13792 ( .A(n8031), .Z(n396) );
  HS65_LS_IVX2 U13793 ( .A(n5393), .Z(n483) );
  HS65_LS_IVX2 U13794 ( .A(n5161), .Z(n701) );
  HS65_LS_IVX2 U13795 ( .A(n5039), .Z(n37) );
  HS65_LS_IVX2 U13796 ( .A(n6985), .Z(n306) );
  HS65_LS_IVX2 U13797 ( .A(n6753), .Z(n519) );
  HS65_LS_IVX2 U13798 ( .A(n6870), .Z(n85) );
  HS65_LS_IVX2 U13799 ( .A(n6632), .Z(n563) );
  HS65_LS_IVX2 U13800 ( .A(n5278), .Z(n264) );
  HS65_LS_IVX2 U13801 ( .A(n2529), .Z(n903) );
  HS65_LS_IVX2 U13802 ( .A(n1777), .Z(n821) );
  HS65_LS_IVX2 U13803 ( .A(n3043), .Z(n172) );
  HS65_LS_IVX2 U13804 ( .A(n8335), .Z(n356) );
  HS65_LS_IVX2 U13805 ( .A(n1401), .Z(n862) );
  HS65_LS_IVX2 U13806 ( .A(n2153), .Z(n780) );
  HS65_LS_NOR2X2 U13807 ( .A(n3064), .B(n3045), .Z(n3664) );
  HS65_LS_IVX2 U13808 ( .A(n7633), .Z(n615) );
  HS65_LS_IVX2 U13809 ( .A(n7661), .Z(n128) );
  HS65_LS_IVX2 U13810 ( .A(n3985), .Z(n438) );
  HS65_LS_IVX2 U13811 ( .A(n3962), .Z(n659) );
  HS65_LS_IVX2 U13812 ( .A(n8542), .Z(n358) );
  HS65_LS_IVX2 U13813 ( .A(n4560), .Z(n11) );
  HS65_LS_IVX2 U13814 ( .A(n6153), .Z(n537) );
  HS65_LS_IVX2 U13815 ( .A(n8361), .Z(n350) );
  HS65_LS_IVX2 U13816 ( .A(n6058), .Z(n70) );
  HS65_LS_IVX2 U13817 ( .A(n6104), .Z(n291) );
  HS65_LS_IVX2 U13818 ( .A(n4511), .Z(n468) );
  HS65_LS_IVX2 U13819 ( .A(n4465), .Z(n249) );
  HS65_LS_IVX2 U13820 ( .A(n4636), .Z(n676) );
  HS65_LS_IVX2 U13821 ( .A(n6229), .Z(n494) );
  HS65_LS_IVX2 U13822 ( .A(n3585), .Z(n177) );
  HS65_LS_IVX2 U13823 ( .A(n8881), .Z(n341) );
  HS65_LS_NOR2X2 U13824 ( .A(n6313), .B(n7108), .Z(n6673) );
  HS65_LS_NOR2X2 U13825 ( .A(n4720), .B(n5516), .Z(n5080) );
  HS65_LS_NOR2X2 U13826 ( .A(n2256), .B(n2528), .Z(n2309) );
  HS65_LS_NOR2X2 U13827 ( .A(n1504), .B(n1776), .Z(n1557) );
  HS65_LS_OAI212X3 U13828 ( .A(n8428), .B(n7793), .C(n7847), .D(n8160), .E(
        n8429), .Z(n8419) );
  HS65_LS_NOR2X2 U13829 ( .A(n594), .B(n597), .Z(n8428) );
  HS65_LS_OAI21X2 U13830 ( .A(n601), .B(n591), .C(n615), .Z(n8429) );
  HS65_LS_OAI212X3 U13831 ( .A(n8488), .B(n7893), .C(n7886), .D(n8192), .E(
        n8489), .Z(n8479) );
  HS65_LS_NOR2X2 U13832 ( .A(n107), .B(n110), .Z(n8488) );
  HS65_LS_OAI21X2 U13833 ( .A(n114), .B(n104), .C(n128), .Z(n8489) );
  HS65_LS_IVX2 U13834 ( .A(n7109), .Z(n569) );
  HS65_LS_IVX2 U13835 ( .A(n5517), .Z(n43) );
  HS65_LS_NAND2X2 U13836 ( .A(n2965), .B(n3905), .Z(n3085) );
  HS65_LS_IVX2 U13837 ( .A(n8070), .Z(n353) );
  HS65_LS_IVX2 U13838 ( .A(n1548), .Z(n844) );
  HS65_LS_IVX2 U13839 ( .A(n2300), .Z(n926) );
  HS65_LS_NOR2X2 U13840 ( .A(n1128), .B(n1400), .Z(n1181) );
  HS65_LS_NOR2X2 U13841 ( .A(n1880), .B(n2152), .Z(n1933) );
  HS65_LS_OAI212X3 U13842 ( .A(n8541), .B(n8542), .C(n8543), .D(n7778), .E(
        n8544), .Z(n8530) );
  HS65_LS_NOR2X2 U13843 ( .A(n330), .B(n326), .Z(n8541) );
  HS65_LS_NAND2X2 U13844 ( .A(n8045), .B(n7953), .Z(n8346) );
  HS65_LS_IVX2 U13845 ( .A(n7793), .Z(n618) );
  HS65_LS_IVX2 U13846 ( .A(n7893), .Z(n131) );
  HS65_LS_IVX2 U13847 ( .A(n3940), .Z(n213) );
  HS65_LS_AOI212X2 U13848 ( .A(n16), .B(n5086), .C(n42), .D(n26), .E(n5726), 
        .Z(n5725) );
  HS65_LS_CBI4I1X3 U13849 ( .A(n4562), .B(n4488), .C(n4577), .D(n5123), .Z(
        n5726) );
  HS65_LS_AOI212X2 U13850 ( .A(n542), .B(n6679), .C(n568), .D(n552), .E(n7318), 
        .Z(n7317) );
  HS65_LS_CBI4I1X3 U13851 ( .A(n6155), .B(n6081), .C(n6170), .D(n6716), .Z(
        n7318) );
  HS65_LS_IVX2 U13852 ( .A(n3964), .Z(n662) );
  HS65_LS_IVX2 U13853 ( .A(n2504), .Z(n897) );
  HS65_LS_IVX2 U13854 ( .A(n1376), .Z(n856) );
  HS65_LS_IVX2 U13855 ( .A(n2128), .Z(n774) );
  HS65_LS_IVX2 U13856 ( .A(n1752), .Z(n815) );
  HS65_LS_IVX2 U13857 ( .A(n3536), .Z(n222) );
  HS65_LS_NOR2X2 U13858 ( .A(n3940), .B(n2965), .Z(n3497) );
  HS65_LS_IVX2 U13859 ( .A(n3942), .Z(n210) );
  HS65_LS_NOR2X2 U13860 ( .A(n2848), .B(n3983), .Z(n3197) );
  HS65_LS_IVX2 U13861 ( .A(n6288), .Z(n568) );
  HS65_LS_IVX2 U13862 ( .A(n4695), .Z(n42) );
  HS65_LS_IVX2 U13863 ( .A(n1686), .Z(n818) );
  HS65_LS_IVX2 U13864 ( .A(n2438), .Z(n900) );
  HS65_LS_NOR2X2 U13865 ( .A(n3264), .B(n3045), .Z(n3665) );
  HS65_LS_IVX2 U13866 ( .A(n2901), .Z(n670) );
  HS65_LS_IVX2 U13867 ( .A(n8095), .Z(n391) );
  HS65_LS_IVX2 U13868 ( .A(n1172), .Z(n885) );
  HS65_LS_IVX2 U13869 ( .A(n1924), .Z(n803) );
  HS65_LS_IVX2 U13870 ( .A(n1310), .Z(n859) );
  HS65_LS_IVX2 U13871 ( .A(n1776), .Z(n822) );
  HS65_LS_IVX2 U13872 ( .A(n2528), .Z(n904) );
  HS65_LS_IVX2 U13873 ( .A(n5523), .Z(n32) );
  HS65_LS_IVX2 U13874 ( .A(n7115), .Z(n558) );
  HS65_LS_IVX2 U13875 ( .A(n3188), .Z(n412) );
  HS65_LS_IVX2 U13876 ( .A(n7646), .Z(n599) );
  HS65_LS_IVX2 U13877 ( .A(n7674), .Z(n112) );
  HS65_LS_IVX2 U13878 ( .A(n2062), .Z(n777) );
  HS65_LS_NOR2X2 U13879 ( .A(n4576), .B(n5516), .Z(n4704) );
  HS65_LS_NOR2X2 U13880 ( .A(n6169), .B(n7108), .Z(n6297) );
  HS65_LS_IVX2 U13881 ( .A(n1400), .Z(n863) );
  HS65_LS_IVX2 U13882 ( .A(n2152), .Z(n781) );
  HS65_LS_IVX2 U13883 ( .A(n3045), .Z(n157) );
  HS65_LS_OAI212X3 U13884 ( .A(n3584), .B(n3585), .C(n3586), .D(n3281), .E(
        n3587), .Z(n3573) );
  HS65_LS_NOR2X2 U13885 ( .A(n156), .B(n159), .Z(n3584) );
  HS65_LS_IVX2 U13886 ( .A(n6339), .Z(n60) );
  HS65_LS_IVX2 U13887 ( .A(n4785), .Z(n458) );
  HS65_LS_IVX2 U13888 ( .A(n6378), .Z(n281) );
  HS65_LS_IVX2 U13889 ( .A(n4746), .Z(n239) );
  HS65_LS_IVX2 U13890 ( .A(n4639), .Z(n683) );
  HS65_LS_IVX2 U13891 ( .A(n6232), .Z(n501) );
  HS65_LS_IVX2 U13892 ( .A(n7663), .Z(n133) );
  HS65_LS_IVX2 U13893 ( .A(n7635), .Z(n620) );
  HS65_LS_IVX2 U13894 ( .A(n2323), .Z(n928) );
  HS65_LS_IVX2 U13895 ( .A(n1571), .Z(n846) );
  HS65_LS_NOR2X2 U13896 ( .A(n8159), .B(n7639), .Z(n8399) );
  HS65_LS_NOR2X2 U13897 ( .A(n8191), .B(n7667), .Z(n8459) );
  HS65_LS_NOR2X2 U13898 ( .A(n3100), .B(n2965), .Z(n3438) );
  HS65_LS_IVX2 U13899 ( .A(n2856), .Z(n446) );
  HS65_LS_IVX2 U13900 ( .A(n3074), .Z(n221) );
  HS65_LS_IVX2 U13901 ( .A(n3983), .Z(n435) );
  HS65_LS_NOR2X2 U13902 ( .A(n8639), .B(n8045), .Z(n8581) );
  HS65_LS_OAI212X3 U13903 ( .A(n3483), .B(n3484), .C(n2875), .D(n2878), .E(
        n3485), .Z(n3473) );
  HS65_LS_NOR2X2 U13904 ( .A(n197), .B(n3426), .Z(n3483) );
  HS65_LS_IVX2 U13905 ( .A(n1195), .Z(n887) );
  HS65_LS_IVX2 U13906 ( .A(n1947), .Z(n805) );
  HS65_LS_IVX2 U13907 ( .A(n5639), .Z(n477) );
  HS65_LS_IVX2 U13908 ( .A(n5612), .Z(n258) );
  HS65_LS_IVX2 U13909 ( .A(n7231), .Z(n300) );
  HS65_LS_IVX2 U13910 ( .A(n7204), .Z(n79) );
  HS65_LS_IVX2 U13911 ( .A(n5588), .Z(n696) );
  HS65_LS_IVX2 U13912 ( .A(n7180), .Z(n514) );
  HS65_LS_IVX2 U13913 ( .A(n2927), .Z(n159) );
  HS65_LS_IVX2 U13914 ( .A(n3280), .Z(n170) );
  HS65_LS_IVX2 U13915 ( .A(n6155), .Z(n544) );
  HS65_LS_IVX2 U13916 ( .A(n4562), .Z(n18) );
  HS65_LS_IVX2 U13917 ( .A(n2972), .Z(n218) );
  HS65_LS_NOR2X2 U13918 ( .A(n4576), .B(n5517), .Z(n4713) );
  HS65_LS_NOR2X2 U13919 ( .A(n6169), .B(n7109), .Z(n6306) );
  HS65_LS_IVX2 U13920 ( .A(n3147), .Z(n635) );
  HS65_LS_IVX2 U13921 ( .A(n2945), .Z(n202) );
  HS65_LS_IVX2 U13922 ( .A(n2943), .Z(n190) );
  HS65_LS_NOR2X2 U13923 ( .A(n7858), .B(n8009), .Z(n8301) );
  HS65_LS_IVX2 U13924 ( .A(n3042), .Z(n144) );
  HS65_LS_IVX2 U13925 ( .A(n8040), .Z(n336) );
  HS65_LS_NOR2X2 U13926 ( .A(n2923), .B(n3264), .Z(n3637) );
  HS65_LS_IVX2 U13927 ( .A(n3203), .Z(n421) );
  HS65_LS_IVX2 U13928 ( .A(n8004), .Z(n374) );
  HS65_LS_NOR2X2 U13929 ( .A(n8160), .B(n7635), .Z(n7809) );
  HS65_LS_NOR2X2 U13930 ( .A(n8192), .B(n7663), .Z(n7909) );
  HS65_LS_AOI212X2 U13931 ( .A(n880), .B(n859), .C(n888), .D(n864), .E(n1120), 
        .Z(n1119) );
  HS65_LS_OAI21X2 U13932 ( .A(n1121), .B(n1122), .C(n1123), .Z(n1120) );
  HS65_LS_AOI212X2 U13933 ( .A(n798), .B(n777), .C(n806), .D(n782), .E(n1872), 
        .Z(n1871) );
  HS65_LS_OAI21X2 U13934 ( .A(n1873), .B(n1874), .C(n1875), .Z(n1872) );
  HS65_LS_IVX2 U13935 ( .A(n8046), .Z(n324) );
  HS65_LS_IVX2 U13936 ( .A(n3064), .Z(n176) );
  HS65_LS_NAND2X2 U13937 ( .A(n4581), .B(n5492), .Z(n4693) );
  HS65_LS_NAND2X2 U13938 ( .A(n6174), .B(n7084), .Z(n6286) );
  HS65_LS_OAI212X3 U13939 ( .A(n8975), .B(n8252), .C(n8031), .D(n8220), .E(
        n8976), .Z(n8974) );
  HS65_LS_OAI21X2 U13940 ( .A(n381), .B(n373), .C(n394), .Z(n8976) );
  HS65_LS_NOR3X1 U13941 ( .A(n397), .B(n388), .C(n390), .Z(n8975) );
  HS65_LS_IVX2 U13942 ( .A(n3236), .Z(n175) );
  HS65_LS_NAND2X2 U13943 ( .A(n6358), .B(n6064), .Z(n6503) );
  HS65_LS_NAND2X2 U13944 ( .A(n6397), .B(n6110), .Z(n6557) );
  HS65_LS_NAND2X2 U13945 ( .A(n4804), .B(n4517), .Z(n4964) );
  HS65_LS_NAND2X2 U13946 ( .A(n4765), .B(n4471), .Z(n4910) );
  HS65_LS_NAND2X2 U13947 ( .A(n4658), .B(n5508), .Z(n4833) );
  HS65_LS_NAND2X2 U13948 ( .A(n6251), .B(n7100), .Z(n6426) );
  HS65_LS_NOR2X2 U13949 ( .A(n3962), .B(n3167), .Z(n3739) );
  HS65_LS_OAI212X3 U13950 ( .A(n1194), .B(n1195), .C(n1196), .D(n1128), .E(
        n1197), .Z(n1190) );
  HS65_LS_AOI12X2 U13951 ( .A(n853), .B(n1198), .C(n1199), .Z(n1197) );
  HS65_LS_AOI12X2 U13952 ( .A(n1200), .B(n1172), .C(n1201), .Z(n1199) );
  HS65_LS_OAI212X3 U13953 ( .A(n1946), .B(n1947), .C(n1948), .D(n1880), .E(
        n1949), .Z(n1942) );
  HS65_LS_AOI12X2 U13954 ( .A(n771), .B(n1950), .C(n1951), .Z(n1949) );
  HS65_LS_AOI12X2 U13955 ( .A(n1952), .B(n1924), .C(n1953), .Z(n1951) );
  HS65_LS_AOI212X2 U13956 ( .A(n656), .B(n3695), .C(n666), .D(n3696), .E(n3697), .Z(n3694) );
  HS65_LS_NAND2X2 U13957 ( .A(n2984), .B(n2893), .Z(n3696) );
  HS65_LS_NAND2X2 U13958 ( .A(n3167), .B(n2900), .Z(n3314) );
  HS65_LS_NAND4ABX3 U13959 ( .A(n2931), .B(n2932), .C(n2933), .D(n2934), .Z(
        n2652) );
  HS65_LS_NAND4ABX3 U13960 ( .A(n2967), .B(n2968), .C(n2969), .D(n2970), .Z(
        n2931) );
  HS65_LS_OAI212X3 U13961 ( .A(n2959), .B(n2960), .C(n2961), .D(n2878), .E(
        n2962), .Z(n2932) );
  HS65_LS_AOI212X2 U13962 ( .A(n189), .B(n215), .C(n193), .D(n212), .E(n2935), 
        .Z(n2934) );
  HS65_LS_IVX2 U13963 ( .A(n3162), .Z(n645) );
  HS65_LS_AOI212X2 U13964 ( .A(n462), .B(n5439), .C(n489), .D(n456), .E(n5903), 
        .Z(n5902) );
  HS65_LS_CBI4I1X3 U13965 ( .A(n4785), .B(n4510), .C(n4800), .D(n5460), .Z(
        n5903) );
  HS65_LS_AOI212X2 U13966 ( .A(n243), .B(n5324), .C(n270), .D(n237), .E(n5844), 
        .Z(n5843) );
  HS65_LS_CBI4I1X3 U13967 ( .A(n4746), .B(n4464), .C(n4761), .D(n5345), .Z(
        n5844) );
  HS65_LS_AOI212X2 U13968 ( .A(n681), .B(n5208), .C(n706), .D(n690), .E(n5788), 
        .Z(n5787) );
  HS65_LS_CBI4I1X3 U13969 ( .A(n4639), .B(n4544), .C(n4654), .D(n5229), .Z(
        n5788) );
  HS65_LS_AOI212X2 U13970 ( .A(n285), .B(n7031), .C(n312), .D(n279), .E(n7495), 
        .Z(n7494) );
  HS65_LS_CBI4I1X3 U13971 ( .A(n6378), .B(n6103), .C(n6393), .D(n7052), .Z(
        n7495) );
  HS65_LS_AOI212X2 U13972 ( .A(n499), .B(n6800), .C(n524), .D(n508), .E(n7380), 
        .Z(n7379) );
  HS65_LS_CBI4I1X3 U13973 ( .A(n6232), .B(n6137), .C(n6247), .D(n6821), .Z(
        n7380) );
  HS65_LS_AOI212X2 U13974 ( .A(n64), .B(n6916), .C(n91), .D(n58), .E(n7436), 
        .Z(n7435) );
  HS65_LS_CBI4I1X3 U13975 ( .A(n6339), .B(n6057), .C(n6354), .D(n6937), .Z(
        n7436) );
  HS65_LS_NOR2X2 U13976 ( .A(n8663), .B(n8003), .Z(n8277) );
  HS65_LS_IVX2 U13977 ( .A(n3052), .Z(n150) );
  HS65_LS_OAI212X3 U13978 ( .A(n1793), .B(n1510), .C(n1686), .D(n1529), .E(
        n1794), .Z(n1792) );
  HS65_LS_NOR3X1 U13979 ( .A(n814), .B(n823), .C(n816), .Z(n1793) );
  HS65_LS_OAI21X2 U13980 ( .A(n839), .B(n846), .C(n828), .Z(n1794) );
  HS65_LS_OAI212X3 U13981 ( .A(n2545), .B(n2262), .C(n2438), .D(n2281), .E(
        n2546), .Z(n2544) );
  HS65_LS_NOR3X1 U13982 ( .A(n896), .B(n905), .C(n898), .Z(n2545) );
  HS65_LS_OAI21X2 U13983 ( .A(n921), .B(n928), .C(n910), .Z(n2546) );
  HS65_LS_IVX2 U13984 ( .A(n7998), .Z(n373) );
  HS65_LS_NAND2X2 U13985 ( .A(n8003), .B(n7870), .Z(n8093) );
  HS65_LS_NOR2X2 U13986 ( .A(n7833), .B(n8160), .Z(n8758) );
  HS65_LS_NOR2X2 U13987 ( .A(n7932), .B(n8192), .Z(n8846) );
  HS65_LS_IVX2 U13988 ( .A(n2895), .Z(n650) );
  HS65_LS_AOI212X2 U13989 ( .A(n96), .B(n7915), .C(n109), .D(n131), .E(n7916), 
        .Z(n7914) );
  HS65_LS_CBI4I1X3 U13990 ( .A(n7674), .B(n7880), .C(n7917), .D(n7918), .Z(
        n7916) );
  HS65_LS_AOI212X2 U13991 ( .A(n583), .B(n7815), .C(n596), .D(n618), .E(n7816), 
        .Z(n7814) );
  HS65_LS_CBI4I1X3 U13992 ( .A(n7646), .B(n7817), .C(n7818), .D(n7819), .Z(
        n7816) );
  HS65_LS_IVX2 U13993 ( .A(n6065), .Z(n88) );
  HS65_LS_IVX2 U13994 ( .A(n4472), .Z(n267) );
  HS65_LS_IVX2 U13995 ( .A(n4518), .Z(n486) );
  HS65_LS_IVX2 U13996 ( .A(n6111), .Z(n309) );
  HS65_LS_IVX2 U13997 ( .A(n6126), .Z(n523) );
  HS65_LS_IVX2 U13998 ( .A(n4533), .Z(n705) );
  HS65_LS_NOR2X2 U13999 ( .A(n3905), .B(n2961), .Z(n3478) );
  HS65_LS_OAI212X3 U14000 ( .A(n1417), .B(n1134), .C(n1310), .D(n1153), .E(
        n1418), .Z(n1416) );
  HS65_LS_NOR3X1 U14001 ( .A(n855), .B(n864), .C(n857), .Z(n1417) );
  HS65_LS_OAI21X2 U14002 ( .A(n880), .B(n887), .C(n869), .Z(n1418) );
  HS65_LS_OAI212X3 U14003 ( .A(n2169), .B(n1886), .C(n2062), .D(n1905), .E(
        n2170), .Z(n2168) );
  HS65_LS_NOR3X1 U14004 ( .A(n773), .B(n782), .C(n775), .Z(n2169) );
  HS65_LS_OAI21X2 U14005 ( .A(n798), .B(n805), .C(n787), .Z(n2170) );
  HS65_LS_NOR2X2 U14006 ( .A(n6353), .B(n7137), .Z(n6513) );
  HS65_LS_NOR2X2 U14007 ( .A(n6392), .B(n7158), .Z(n6567) );
  HS65_LS_NOR2X2 U14008 ( .A(n4799), .B(n5566), .Z(n4974) );
  HS65_LS_NOR2X2 U14009 ( .A(n4760), .B(n5545), .Z(n4920) );
  HS65_LS_NOR2X2 U14010 ( .A(n4653), .B(n5581), .Z(n4844) );
  HS65_LS_NOR2X2 U14011 ( .A(n6246), .B(n7173), .Z(n6437) );
  HS65_LS_IVX2 U14012 ( .A(n6086), .Z(n567) );
  HS65_LS_IVX2 U14013 ( .A(n4493), .Z(n41) );
  HS65_LS_IVX2 U14014 ( .A(n8160), .Z(n586) );
  HS65_LS_IVX2 U14015 ( .A(n8192), .Z(n99) );
  HS65_LS_IVX2 U14016 ( .A(n8009), .Z(n399) );
  HS65_LS_NOR2X2 U14017 ( .A(n2894), .B(n3167), .Z(n3682) );
  HS65_LS_OAI212X3 U14018 ( .A(n4040), .B(n2854), .C(n3843), .D(n3002), .E(
        n4041), .Z(n4039) );
  HS65_LS_NOR3X1 U14019 ( .A(n442), .B(n434), .C(n430), .Z(n4040) );
  HS65_LS_OAI21X2 U14020 ( .A(n417), .B(n421), .C(n446), .Z(n4041) );
  HS65_LS_OAI212X3 U14021 ( .A(n7930), .B(n7662), .C(n7931), .D(n7932), .E(
        n7933), .Z(n7929) );
  HS65_LS_NOR3X1 U14022 ( .A(n119), .B(n125), .C(n124), .Z(n7930) );
  HS65_LS_OAI21X2 U14023 ( .A(n106), .B(n99), .C(n132), .Z(n7933) );
  HS65_LS_OAI212X3 U14024 ( .A(n8915), .B(n8556), .C(n8070), .D(n8525), .E(
        n8916), .Z(n8914) );
  HS65_LS_OAI21X2 U14025 ( .A(n332), .B(n336), .C(n356), .Z(n8916) );
  HS65_LS_NOR3X1 U14026 ( .A(n350), .B(n348), .C(n349), .Z(n8915) );
  HS65_LS_NOR2X2 U14027 ( .A(n2924), .B(n3064), .Z(n3568) );
  HS65_LS_NOR2X2 U14028 ( .A(n3536), .B(n2960), .Z(n3099) );
  HS65_LS_NOR2X2 U14029 ( .A(n3236), .B(n3042), .Z(n3261) );
  HS65_LS_NAND4ABX3 U14030 ( .A(n3068), .B(n3069), .C(n3070), .D(n3071), .Z(
        n2740) );
  HS65_LS_OAI212X3 U14031 ( .A(n3125), .B(n2943), .C(n3126), .D(n3127), .E(
        n3128), .Z(n3069) );
  HS65_LS_NAND4ABX3 U14032 ( .A(n3129), .B(n3130), .C(n3131), .D(n3132), .Z(
        n3068) );
  HS65_LS_AOI212X2 U14033 ( .A(n203), .B(n3072), .C(n228), .D(n198), .E(n3073), 
        .Z(n3071) );
  HS65_LS_NAND4ABX3 U14034 ( .A(n8493), .B(n8494), .C(n8495), .D(n8496), .Z(
        n2763) );
  HS65_LS_CB4I6X4 U14035 ( .A(n401), .B(n397), .C(n381), .D(n8286), .Z(n8493)
         );
  HS65_LS_AOI212X2 U14036 ( .A(n374), .B(n398), .C(n376), .D(n8506), .E(n8507), 
        .Z(n8495) );
  HS65_LS_CBI4I1X3 U14037 ( .A(n389), .B(n7762), .C(n7861), .D(n8508), .Z(
        n8494) );
  HS65_LS_OAI212X3 U14038 ( .A(n4016), .B(n2899), .C(n3726), .D(n2984), .E(
        n4017), .Z(n4015) );
  HS65_LS_OAI21X2 U14039 ( .A(n641), .B(n645), .C(n670), .Z(n4017) );
  HS65_LS_NOR3X1 U14040 ( .A(n666), .B(n658), .C(n654), .Z(n4016) );
  HS65_LS_NOR2X2 U14041 ( .A(n7953), .B(n8041), .Z(n8564) );
  HS65_LS_NOR2X2 U14042 ( .A(n3776), .B(n3162), .Z(n3327) );
  HS65_LS_OAI212X3 U14043 ( .A(n5632), .B(n4516), .C(n4620), .D(n5393), .E(
        n5633), .Z(n5631) );
  HS65_LS_NOR3X1 U14044 ( .A(n484), .B(n471), .C(n475), .Z(n5632) );
  HS65_LS_OAI21X2 U14045 ( .A(n455), .B(n463), .C(n486), .Z(n5633) );
  HS65_LS_OAI212X3 U14046 ( .A(n5605), .B(n4470), .C(n4595), .D(n5278), .E(
        n5606), .Z(n5604) );
  HS65_LS_NOR3X1 U14047 ( .A(n265), .B(n252), .C(n256), .Z(n5605) );
  HS65_LS_OAI21X2 U14048 ( .A(n236), .B(n244), .C(n267), .Z(n5606) );
  HS65_LS_OAI212X3 U14049 ( .A(n7224), .B(n6109), .C(n6213), .D(n6985), .E(
        n7225), .Z(n7223) );
  HS65_LS_NOR3X1 U14050 ( .A(n307), .B(n294), .C(n298), .Z(n7224) );
  HS65_LS_OAI21X2 U14051 ( .A(n278), .B(n286), .C(n309), .Z(n7225) );
  HS65_LS_OAI212X3 U14052 ( .A(n5781), .B(n4535), .C(n5148), .D(n5161), .E(
        n5782), .Z(n5780) );
  HS65_LS_NOR3X1 U14053 ( .A(n699), .B(n711), .C(n709), .Z(n5781) );
  HS65_LS_OAI21X2 U14054 ( .A(n689), .B(n682), .C(n705), .Z(n5782) );
  HS65_LS_OAI212X3 U14055 ( .A(n5719), .B(n4495), .C(n5026), .D(n5039), .E(
        n5720), .Z(n5718) );
  HS65_LS_OAI21X2 U14056 ( .A(n25), .B(n17), .C(n41), .Z(n5720) );
  HS65_LS_NOR3X1 U14057 ( .A(n45), .B(n47), .C(n35), .Z(n5719) );
  HS65_LS_OAI212X3 U14058 ( .A(n7373), .B(n6128), .C(n6740), .D(n6753), .E(
        n7374), .Z(n7372) );
  HS65_LS_NOR3X1 U14059 ( .A(n517), .B(n529), .C(n527), .Z(n7373) );
  HS65_LS_OAI21X2 U14060 ( .A(n507), .B(n500), .C(n523), .Z(n7374) );
  HS65_LS_OAI212X3 U14061 ( .A(n7197), .B(n6063), .C(n6188), .D(n6870), .E(
        n7198), .Z(n7196) );
  HS65_LS_NOR3X1 U14062 ( .A(n86), .B(n73), .C(n77), .Z(n7197) );
  HS65_LS_OAI21X2 U14063 ( .A(n57), .B(n65), .C(n88), .Z(n7198) );
  HS65_LS_OAI212X3 U14064 ( .A(n7311), .B(n6088), .C(n6619), .D(n6632), .E(
        n7312), .Z(n7310) );
  HS65_LS_OAI21X2 U14065 ( .A(n551), .B(n543), .C(n567), .Z(n7312) );
  HS65_LS_NOR3X1 U14066 ( .A(n571), .B(n573), .C(n561), .Z(n7311) );
  HS65_LS_IVX2 U14067 ( .A(n2960), .Z(n195) );
  HS65_LS_NOR2X2 U14068 ( .A(n8412), .B(n7793), .Z(n8757) );
  HS65_LS_NOR2X2 U14069 ( .A(n8472), .B(n7893), .Z(n8845) );
  HS65_LS_IVX2 U14070 ( .A(n4576), .Z(n17) );
  HS65_LS_IVX2 U14071 ( .A(n6169), .Z(n543) );
  HS65_LS_IVX2 U14072 ( .A(n4581), .Z(n16) );
  HS65_LS_IVX2 U14073 ( .A(n6174), .Z(n542) );
  HS65_LS_IVX2 U14074 ( .A(n4653), .Z(n682) );
  HS65_LS_IVX2 U14075 ( .A(n4799), .Z(n463) );
  HS65_LS_IVX2 U14076 ( .A(n6392), .Z(n286) );
  HS65_LS_IVX2 U14077 ( .A(n6353), .Z(n65) );
  HS65_LS_IVX2 U14078 ( .A(n6246), .Z(n500) );
  HS65_LS_IVX2 U14079 ( .A(n4760), .Z(n244) );
  HS65_LS_IVX2 U14080 ( .A(n3215), .Z(n439) );
  HS65_LS_NOR2X2 U14081 ( .A(n2263), .B(n2324), .Z(n2432) );
  HS65_LS_NOR2X2 U14082 ( .A(n1511), .B(n1572), .Z(n1680) );
  HS65_LS_NAND2X2 U14083 ( .A(n6056), .B(n6050), .Z(n6489) );
  HS65_LS_NAND2X2 U14084 ( .A(n6102), .B(n6096), .Z(n6543) );
  HS65_LS_NAND2X2 U14085 ( .A(n4463), .B(n4457), .Z(n4896) );
  HS65_LS_NAND2X2 U14086 ( .A(n4509), .B(n4503), .Z(n4950) );
  HS65_LS_NAND2X2 U14087 ( .A(n4862), .B(n4835), .Z(n4818) );
  HS65_LS_NAND2X2 U14088 ( .A(n6455), .B(n6428), .Z(n6411) );
  HS65_LS_NOR2X2 U14089 ( .A(n7870), .B(n7999), .Z(n8260) );
  HS65_LS_NOR2X2 U14090 ( .A(n1135), .B(n1196), .Z(n1304) );
  HS65_LS_NOR2X2 U14091 ( .A(n1887), .B(n1948), .Z(n2056) );
  HS65_LS_NOR2X2 U14092 ( .A(n2887), .B(n3147), .Z(n3759) );
  HS65_LS_NOR2X2 U14093 ( .A(n4799), .B(n5393), .Z(n5471) );
  HS65_LS_NOR2X2 U14094 ( .A(n4760), .B(n5278), .Z(n5356) );
  HS65_LS_NOR2X2 U14095 ( .A(n6392), .B(n6985), .Z(n7063) );
  HS65_LS_NOR2X2 U14096 ( .A(n4653), .B(n5161), .Z(n5241) );
  HS65_LS_NOR2X2 U14097 ( .A(n4576), .B(n5039), .Z(n5105) );
  HS65_LS_NOR2X2 U14098 ( .A(n6246), .B(n6753), .Z(n6833) );
  HS65_LS_NOR2X2 U14099 ( .A(n6353), .B(n6870), .Z(n6948) );
  HS65_LS_NOR2X2 U14100 ( .A(n6169), .B(n6632), .Z(n6698) );
  HS65_LS_NAND4ABX3 U14101 ( .A(n8074), .B(n8075), .C(n8076), .D(n8077), .Z(
        n2765) );
  HS65_LS_OAI212X3 U14102 ( .A(n8129), .B(n7872), .C(n368), .D(n8130), .E(
        n8131), .Z(n8075) );
  HS65_LS_NAND4ABX3 U14103 ( .A(n8132), .B(n8133), .C(n8134), .D(n8135), .Z(
        n8074) );
  HS65_LS_AOI212X2 U14104 ( .A(n376), .B(n8078), .C(n380), .D(n386), .E(n8079), 
        .Z(n8077) );
  HS65_LS_NOR2X2 U14105 ( .A(n2855), .B(n3204), .Z(n3837) );
  HS65_LS_NOR2X2 U14106 ( .A(n7881), .B(n8192), .Z(n7935) );
  HS65_LS_NOR2X2 U14107 ( .A(n7842), .B(n8160), .Z(n7836) );
  HS65_LS_IVX2 U14108 ( .A(n4804), .Z(n462) );
  HS65_LS_IVX2 U14109 ( .A(n4765), .Z(n243) );
  HS65_LS_IVX2 U14110 ( .A(n4658), .Z(n681) );
  HS65_LS_IVX2 U14111 ( .A(n6397), .Z(n285) );
  HS65_LS_IVX2 U14112 ( .A(n6358), .Z(n64) );
  HS65_LS_IVX2 U14113 ( .A(n6251), .Z(n499) );
  HS65_LS_NOR2AX3 U14114 ( .A(n7709), .B(n8150), .Z(n7708) );
  HS65_LS_NOR2AX3 U14115 ( .A(n7747), .B(n8182), .Z(n7746) );
  HS65_LS_NOR2X2 U14116 ( .A(n2900), .B(n3163), .Z(n3721) );
  HS65_LS_NAND4ABX3 U14117 ( .A(n4006), .B(n4007), .C(n4008), .D(n4009), .Z(
        n2757) );
  HS65_LS_CB4I6X4 U14118 ( .A(n660), .B(n659), .C(n635), .D(n3743), .Z(n4006)
         );
  HS65_LS_AOI222X2 U14119 ( .A(n646), .B(n666), .C(n633), .D(n4028), .E(n639), 
        .F(n662), .Z(n4008) );
  HS65_LS_CBI4I1X3 U14120 ( .A(n2990), .B(n3173), .C(n3778), .D(n4029), .Z(
        n4007) );
  HS65_LS_IVX2 U14121 ( .A(n4800), .Z(n475) );
  HS65_LS_IVX2 U14122 ( .A(n4761), .Z(n256) );
  HS65_LS_IVX2 U14123 ( .A(n6393), .Z(n298) );
  HS65_LS_IVX2 U14124 ( .A(n4654), .Z(n709) );
  HS65_LS_IVX2 U14125 ( .A(n6247), .Z(n527) );
  HS65_LS_IVX2 U14126 ( .A(n6354), .Z(n77) );
  HS65_LS_NAND2X2 U14127 ( .A(n3264), .B(n3064), .Z(n3234) );
  HS65_LS_OAI212X3 U14128 ( .A(n3122), .B(n3123), .C(n2960), .D(n3074), .E(
        n3124), .Z(n3112) );
  HS65_LS_OAI21X2 U14129 ( .A(n205), .B(n189), .C(n218), .Z(n3124) );
  HS65_LS_NOR2X2 U14130 ( .A(n199), .B(n198), .Z(n3122) );
  HS65_LS_OAI212X3 U14131 ( .A(n3411), .B(n2842), .C(n3203), .D(n2856), .E(
        n3412), .Z(n3401) );
  HS65_LS_NOR2X2 U14132 ( .A(n415), .B(n414), .Z(n3411) );
  HS65_LS_OAI21X2 U14133 ( .A(n411), .B(n424), .C(n439), .Z(n3412) );
  HS65_LS_NOR2X2 U14134 ( .A(n2923), .B(n4103), .Z(n3618) );
  HS65_LS_NOR2X2 U14135 ( .A(n8315), .B(n7998), .Z(n8118) );
  HS65_LS_NOR2X2 U14136 ( .A(n8159), .B(n7818), .Z(n8762) );
  HS65_LS_NOR2X2 U14137 ( .A(n8191), .B(n7917), .Z(n8850) );
  HS65_LS_NOR2X2 U14138 ( .A(n2875), .B(n2965), .Z(n3526) );
  HS65_LS_NAND4ABX3 U14139 ( .A(n6180), .B(n6181), .C(n6182), .D(n6183), .Z(
        n2799) );
  HS65_LS_CBI4I6X2 U14140 ( .A(n57), .B(n6184), .C(n82), .D(n6185), .Z(n6183)
         );
  HS65_LS_CBI4I1X3 U14141 ( .A(n6194), .B(n6057), .C(n6195), .D(n6196), .Z(
        n6180) );
  HS65_LS_AOI212X2 U14142 ( .A(n76), .B(n65), .C(n91), .D(n58), .E(n6187), .Z(
        n6182) );
  HS65_LS_NAND4ABX3 U14143 ( .A(n4587), .B(n4588), .C(n4589), .D(n4590), .Z(
        n2807) );
  HS65_LS_CBI4I6X2 U14144 ( .A(n236), .B(n4591), .C(n261), .D(n4592), .Z(n4590) );
  HS65_LS_CBI4I1X3 U14145 ( .A(n4601), .B(n4464), .C(n4602), .D(n4603), .Z(
        n4587) );
  HS65_LS_AOI212X2 U14146 ( .A(n255), .B(n244), .C(n270), .D(n237), .E(n4594), 
        .Z(n4589) );
  HS65_LS_IVX2 U14147 ( .A(n8041), .Z(n348) );
  HS65_LS_NOR2X2 U14148 ( .A(n8040), .B(n8361), .Z(n8608) );
  HS65_LS_NOR2X2 U14149 ( .A(n8069), .B(n8070), .Z(n7774) );
  HS65_LS_NAND4ABX3 U14150 ( .A(n2862), .B(n2863), .C(n2864), .D(n2865), .Z(
        n2645) );
  HS65_LS_CBI4I1X3 U14151 ( .A(n2877), .B(n2878), .C(n2879), .D(n2880), .Z(
        n2862) );
  HS65_LS_AOI212X2 U14152 ( .A(n195), .B(n226), .C(n201), .D(n223), .E(n2871), 
        .Z(n2864) );
  HS65_LS_CBI4I1X3 U14153 ( .A(n2873), .B(n2874), .C(n2875), .D(n2876), .Z(
        n2863) );
  HS65_LS_NOR2X2 U14154 ( .A(n2250), .B(n2300), .Z(n2471) );
  HS65_LS_NOR2X2 U14155 ( .A(n1498), .B(n1548), .Z(n1719) );
  HS65_LS_NOR2AX3 U14156 ( .A(n6184), .B(n7204), .Z(n6865) );
  HS65_LS_NOR2AX3 U14157 ( .A(n4616), .B(n5639), .Z(n5388) );
  HS65_LS_NOR2AX3 U14158 ( .A(n4531), .B(n5588), .Z(n5156) );
  HS65_LS_NOR2AX3 U14159 ( .A(n6209), .B(n7231), .Z(n6980) );
  HS65_LS_NOR2AX3 U14160 ( .A(n4591), .B(n5612), .Z(n5273) );
  HS65_LS_NOR2AX3 U14161 ( .A(n6124), .B(n7180), .Z(n6748) );
  HS65_LS_NOR2X2 U14162 ( .A(n4512), .B(n4799), .Z(n5433) );
  HS65_LS_NOR2X2 U14163 ( .A(n4466), .B(n4760), .Z(n5318) );
  HS65_LS_NOR2X2 U14164 ( .A(n6105), .B(n6392), .Z(n7025) );
  HS65_LS_NOR2X2 U14165 ( .A(n4860), .B(n4653), .Z(n5202) );
  HS65_LS_NOR2X2 U14166 ( .A(n6453), .B(n6246), .Z(n6794) );
  HS65_LS_NOR2X2 U14167 ( .A(n6059), .B(n6353), .Z(n6910) );
  HS65_LS_IVX2 U14168 ( .A(n3167), .Z(n644) );
  HS65_LS_NOR2X2 U14169 ( .A(n1122), .B(n1172), .Z(n1343) );
  HS65_LS_NOR2X2 U14170 ( .A(n1874), .B(n1924), .Z(n2095) );
  HS65_LS_NOR2X2 U14171 ( .A(n3065), .B(n2927), .Z(n3620) );
  HS65_LS_IVX2 U14172 ( .A(n8003), .Z(n371) );
  HS65_LS_NAND2X2 U14173 ( .A(n7762), .B(n8095), .Z(n8078) );
  HS65_LS_NAND4ABX3 U14174 ( .A(n7186), .B(n7187), .C(n7188), .D(n7189), .Z(
        n2794) );
  HS65_LS_CB4I6X4 U14175 ( .A(n80), .B(n79), .C(n60), .D(n6893), .Z(n7186) );
  HS65_LS_CBI4I1X3 U14176 ( .A(n6195), .B(n7136), .C(n7210), .D(n7212), .Z(
        n7187) );
  HS65_LS_AOI222X2 U14177 ( .A(n86), .B(n66), .C(n59), .D(n7211), .E(n81), .F(
        n56), .Z(n7188) );
  HS65_LS_NOR2X2 U14178 ( .A(n7857), .B(n8080), .Z(n8124) );
  HS65_LS_NOR2X2 U14179 ( .A(n2842), .B(n3188), .Z(n3876) );
  HS65_LS_IVX2 U14180 ( .A(n3163), .Z(n658) );
  HS65_LS_IVX2 U14181 ( .A(n4577), .Z(n45) );
  HS65_LS_IVX2 U14182 ( .A(n6170), .Z(n571) );
  HS65_LS_NAND4ABX3 U14183 ( .A(n3990), .B(n3991), .C(n3992), .D(n3993), .Z(
        n2907) );
  HS65_LS_CBI4I1X3 U14184 ( .A(n3058), .B(n4002), .C(n3045), .D(n3643), .Z(
        n3990) );
  HS65_LS_CBI4I1X3 U14185 ( .A(n2929), .B(n3065), .C(n3281), .D(n4005), .Z(
        n3991) );
  HS65_LS_AOI222X2 U14186 ( .A(n149), .B(n169), .C(n158), .D(n4004), .E(n154), 
        .F(n165), .Z(n3992) );
  HS65_LS_NOR2X2 U14187 ( .A(n4510), .B(n5639), .Z(n4792) );
  HS65_LS_NOR2X2 U14188 ( .A(n4464), .B(n5612), .Z(n4753) );
  HS65_LS_NOR2X2 U14189 ( .A(n6103), .B(n7231), .Z(n6385) );
  HS65_LS_NOR2X2 U14190 ( .A(n4544), .B(n5588), .Z(n4646) );
  HS65_LS_NOR2X2 U14191 ( .A(n6137), .B(n7180), .Z(n6239) );
  HS65_LS_NOR2X2 U14192 ( .A(n6057), .B(n7204), .Z(n6346) );
  HS65_LS_IVX2 U14193 ( .A(n7999), .Z(n388) );
  HS65_LS_IVX2 U14194 ( .A(n2965), .Z(n197) );
  HS65_LS_IVX2 U14195 ( .A(n2324), .Z(n905) );
  HS65_LS_IVX2 U14196 ( .A(n1572), .Z(n823) );
  HS65_LS_IVX2 U14197 ( .A(n8045), .Z(n337) );
  HS65_LS_IVX2 U14198 ( .A(n1196), .Z(n864) );
  HS65_LS_IVX2 U14199 ( .A(n1948), .Z(n782) );
  HS65_LS_NOR2X2 U14200 ( .A(n3067), .B(n4103), .Z(n3257) );
  HS65_LS_NAND4ABX3 U14201 ( .A(n2974), .B(n2975), .C(n2976), .D(n2977), .Z(
        n2736) );
  HS65_LS_CBI4I1X3 U14202 ( .A(n2985), .B(n2986), .C(n2987), .D(n2988), .Z(
        n2975) );
  HS65_LS_CBI4I1X3 U14203 ( .A(n2989), .B(n2893), .C(n2990), .D(n2991), .Z(
        n2974) );
  HS65_LS_AOI212X2 U14204 ( .A(n645), .B(n656), .C(n640), .D(n669), .E(n2983), 
        .Z(n2976) );
  HS65_LS_NOR2X2 U14205 ( .A(n2923), .B(n3058), .Z(n3256) );
  HS65_LS_IVX2 U14206 ( .A(n3204), .Z(n434) );
  HS65_LS_NAND2X2 U14207 ( .A(n3102), .B(n3123), .Z(n3072) );
  HS65_LS_IVX2 U14208 ( .A(n2985), .Z(n647) );
  HS65_LS_NOR2X2 U14209 ( .A(n3123), .B(n2945), .Z(n3518) );
  HS65_LS_NOR2X2 U14210 ( .A(n1128), .B(n1201), .Z(n1281) );
  HS65_LS_NOR2X2 U14211 ( .A(n2256), .B(n2329), .Z(n2409) );
  HS65_LS_NOR2X2 U14212 ( .A(n1880), .B(n1953), .Z(n2033) );
  HS65_LS_NOR2X2 U14213 ( .A(n1504), .B(n1577), .Z(n1657) );
  HS65_LS_NOR2X2 U14214 ( .A(n6170), .B(n7084), .Z(n6629) );
  HS65_LS_NOR2X2 U14215 ( .A(n4577), .B(n5492), .Z(n5036) );
  HS65_LS_NAND2X2 U14216 ( .A(n3536), .B(n2875), .Z(n3106) );
  HS65_LS_IVX2 U14217 ( .A(n1530), .Z(n837) );
  HS65_LS_IVX2 U14218 ( .A(n2282), .Z(n919) );
  HS65_LS_NAND2X2 U14219 ( .A(n2504), .B(n2284), .Z(n2375) );
  HS65_LS_NAND2X2 U14220 ( .A(n1376), .B(n1156), .Z(n1247) );
  HS65_LS_NAND2X2 U14221 ( .A(n2128), .B(n1908), .Z(n1999) );
  HS65_LS_NAND2X2 U14222 ( .A(n1752), .B(n1532), .Z(n1623) );
  HS65_LS_NOR2X2 U14223 ( .A(n2987), .B(n3167), .Z(n3767) );
  HS65_LS_IVX2 U14224 ( .A(n8164), .Z(n583) );
  HS65_LS_IVX2 U14225 ( .A(n8196), .Z(n96) );
  HS65_LS_IVX2 U14226 ( .A(n1906), .Z(n796) );
  HS65_LS_IVX2 U14227 ( .A(n1154), .Z(n878) );
  HS65_LS_NOR2X2 U14228 ( .A(n3100), .B(n2960), .Z(n3525) );
  HS65_LS_NOR2X2 U14229 ( .A(n2971), .B(n2960), .Z(n3429) );
  HS65_LS_NAND2X2 U14230 ( .A(n7109), .B(n6270), .Z(n6319) );
  HS65_LS_NAND2X2 U14231 ( .A(n5517), .B(n4677), .Z(n4726) );
  HS65_LS_NOR2X2 U14232 ( .A(n1776), .B(n1576), .Z(n1699) );
  HS65_LS_NOR2X2 U14233 ( .A(n2528), .B(n2328), .Z(n2451) );
  HS65_LS_IVX2 U14234 ( .A(n2873), .Z(n192) );
  HS65_LS_NOR2X2 U14235 ( .A(n2152), .B(n1952), .Z(n2075) );
  HS65_LS_NOR2X2 U14236 ( .A(n1400), .B(n1200), .Z(n1323) );
  HS65_LS_NOR2X2 U14237 ( .A(n3983), .B(n3208), .Z(n3856) );
  HS65_LS_NOR2X2 U14238 ( .A(n3063), .B(n3065), .Z(n3636) );
  HS65_LS_NOR2X2 U14239 ( .A(n8030), .B(n8031), .Z(n7757) );
  HS65_LS_NOR2X2 U14240 ( .A(n2856), .B(n3421), .Z(n3880) );
  HS65_LS_NOR2X2 U14241 ( .A(n3074), .B(n3133), .Z(n3522) );
  HS65_LS_OAI212X3 U14242 ( .A(n8700), .B(n7833), .C(n8436), .D(n7817), .E(
        n8701), .Z(n8692) );
  HS65_LS_NOR2X2 U14243 ( .A(n583), .B(n8680), .Z(n8700) );
  HS65_LS_OAI212X3 U14244 ( .A(n8788), .B(n7932), .C(n8447), .D(n7880), .E(
        n8789), .Z(n8780) );
  HS65_LS_NOR2X2 U14245 ( .A(n96), .B(n8768), .Z(n8788) );
  HS65_LS_NOR2X2 U14246 ( .A(n2264), .B(n2281), .Z(n2453) );
  HS65_LS_NOR2X2 U14247 ( .A(n1512), .B(n1529), .Z(n1701) );
  HS65_LS_IVX2 U14248 ( .A(n7917), .Z(n119) );
  HS65_LS_IVX2 U14249 ( .A(n7818), .Z(n606) );
  HS65_LS_IVX2 U14250 ( .A(n3003), .Z(n423) );
  HS65_LS_IVX2 U14251 ( .A(n2961), .Z(n225) );
  HS65_LS_NAND2X2 U14252 ( .A(n7663), .B(n8447), .Z(n7940) );
  HS65_LS_NAND2X2 U14253 ( .A(n7635), .B(n8436), .Z(n7841) );
  HS65_LS_NOR2X2 U14254 ( .A(n1888), .B(n1905), .Z(n2077) );
  HS65_LS_NOR2X2 U14255 ( .A(n1136), .B(n1153), .Z(n1325) );
  HS65_LS_NOR2X2 U14256 ( .A(n4488), .B(n5523), .Z(n4569) );
  HS65_LS_NOR2X2 U14257 ( .A(n6081), .B(n7115), .Z(n6162) );
  HS65_LS_NAND2X2 U14258 ( .A(n7687), .B(n7793), .Z(n8388) );
  HS65_LS_NAND2X2 U14259 ( .A(n7725), .B(n7893), .Z(n8448) );
  HS65_LS_NOR2X2 U14260 ( .A(n2923), .B(n4002), .Z(n3619) );
  HS65_LS_NOR2AX3 U14261 ( .A(n7709), .B(n7793), .Z(n8423) );
  HS65_LS_NOR2AX3 U14262 ( .A(n7747), .B(n7893), .Z(n8483) );
  HS65_LS_NOR2X2 U14263 ( .A(n2945), .B(n2971), .Z(n3521) );
  HS65_LS_NOR2X2 U14264 ( .A(n7778), .B(n8542), .Z(n8524) );
  HS65_LS_NOR2X2 U14265 ( .A(n3074), .B(n3454), .Z(n3500) );
  HS65_LS_NOR2X2 U14266 ( .A(n2856), .B(n3002), .Z(n3858) );
  HS65_LS_NOR2X2 U14267 ( .A(n2901), .B(n2984), .Z(n3741) );
  HS65_LS_NAND2X2 U14268 ( .A(n7191), .B(n6488), .Z(n6533) );
  HS65_LS_NAND2X2 U14269 ( .A(n5599), .B(n4895), .Z(n4940) );
  HS65_LS_NAND2X2 U14270 ( .A(n5626), .B(n5009), .Z(n4994) );
  HS65_LS_NAND2X2 U14271 ( .A(n7218), .B(n6602), .Z(n6587) );
  HS65_LS_NAND2X2 U14272 ( .A(n7174), .B(n6474), .Z(n6459) );
  HS65_LS_NAND2X2 U14273 ( .A(n5582), .B(n4881), .Z(n4866) );
  HS65_LS_IVX2 U14274 ( .A(n8182), .Z(n124) );
  HS65_LS_IVX2 U14275 ( .A(n8150), .Z(n611) );
  HS65_LS_NOR2X2 U14276 ( .A(n7662), .B(n7672), .Z(n7936) );
  HS65_LS_NOR2X2 U14277 ( .A(n7634), .B(n7644), .Z(n7837) );
  HS65_LS_NOR2X2 U14278 ( .A(n8080), .B(n8220), .Z(n7756) );
  HS65_LS_NOR2X2 U14279 ( .A(n2894), .B(n3162), .Z(n3766) );
  HS65_LS_NOR2X2 U14280 ( .A(n8095), .B(n7858), .Z(n8235) );
  HS65_LS_NOR2X2 U14281 ( .A(n2842), .B(n3004), .Z(n3798) );
  HS65_LS_NOR2X2 U14282 ( .A(n7646), .B(n7793), .Z(n8728) );
  HS65_LS_NOR2X2 U14283 ( .A(n7674), .B(n7893), .Z(n8816) );
  HS65_LS_NOR2X2 U14284 ( .A(n6353), .B(n7191), .Z(n6522) );
  HS65_LS_NOR2X2 U14285 ( .A(n6392), .B(n7218), .Z(n6576) );
  HS65_LS_NOR2X2 U14286 ( .A(n4799), .B(n5626), .Z(n4983) );
  HS65_LS_NOR2X2 U14287 ( .A(n4760), .B(n5599), .Z(n4929) );
  HS65_LS_NOR2X2 U14288 ( .A(n4653), .B(n5582), .Z(n4853) );
  HS65_LS_NOR2X2 U14289 ( .A(n6246), .B(n7174), .Z(n6446) );
  HS65_LS_NOR2X2 U14290 ( .A(n6064), .B(n7136), .Z(n6883) );
  HS65_LS_NOR2X2 U14291 ( .A(n4471), .B(n5544), .Z(n5291) );
  HS65_LS_NOR2X2 U14292 ( .A(n4517), .B(n5565), .Z(n5406) );
  HS65_LS_NOR2X2 U14293 ( .A(n6110), .B(n7157), .Z(n6998) );
  HS65_LS_NOR2X2 U14294 ( .A(n5508), .B(n5589), .Z(n5174) );
  HS65_LS_NOR2X2 U14295 ( .A(n7100), .B(n7181), .Z(n6766) );
  HS65_LS_NAND2X2 U14296 ( .A(n4722), .B(n4695), .Z(n4678) );
  HS65_LS_NAND2X2 U14297 ( .A(n6315), .B(n6288), .Z(n6271) );
  HS65_LS_NOR2X2 U14298 ( .A(n2887), .B(n2986), .Z(n3681) );
  HS65_LS_NOR2X2 U14299 ( .A(n3188), .B(n3214), .Z(n3879) );
  HS65_LS_NAND2X2 U14300 ( .A(n2847), .B(n2842), .Z(n3364) );
  HS65_LS_NOR2X2 U14301 ( .A(n8004), .B(n8095), .Z(n8297) );
  HS65_LS_NOR2X2 U14302 ( .A(n7963), .B(n8361), .Z(n8590) );
  HS65_LS_IVX2 U14303 ( .A(n2923), .Z(n147) );
  HS65_LS_NAND2X2 U14304 ( .A(n2892), .B(n2887), .Z(n3302) );
  HS65_LS_NOR2X2 U14305 ( .A(n2440), .B(n2336), .Z(n2354) );
  HS65_LS_NOR2X2 U14306 ( .A(n1688), .B(n1584), .Z(n1602) );
  HS65_LS_NOR2X2 U14307 ( .A(n3123), .B(n2874), .Z(n3437) );
  HS65_LS_NOR2X2 U14308 ( .A(n7084), .B(n7116), .Z(n6645) );
  HS65_LS_NOR2X2 U14309 ( .A(n5492), .B(n5524), .Z(n5052) );
  HS65_LS_AOI212X2 U14310 ( .A(n825), .B(n844), .C(n833), .D(n1517), .E(n1779), 
        .Z(n1760) );
  HS65_LS_AOI12X2 U14311 ( .A(n1497), .B(n1688), .C(n1686), .Z(n1779) );
  HS65_LS_AOI212X2 U14312 ( .A(n907), .B(n926), .C(n915), .D(n2269), .E(n2531), 
        .Z(n2512) );
  HS65_LS_AOI12X2 U14313 ( .A(n2249), .B(n2440), .C(n2438), .Z(n2531) );
  HS65_LS_NOR2X2 U14314 ( .A(n3942), .B(n3101), .Z(n3094) );
  HS65_LS_AOI212X2 U14315 ( .A(n784), .B(n803), .C(n792), .D(n1893), .E(n2155), 
        .Z(n2136) );
  HS65_LS_AOI12X2 U14316 ( .A(n1873), .B(n2064), .C(n2062), .Z(n2155) );
  HS65_LS_AOI212X2 U14317 ( .A(n866), .B(n885), .C(n874), .D(n1141), .E(n1403), 
        .Z(n1384) );
  HS65_LS_AOI12X2 U14318 ( .A(n1121), .B(n1312), .C(n1310), .Z(n1403) );
  HS65_LS_NOR2X2 U14319 ( .A(n4582), .B(n4676), .Z(n5033) );
  HS65_LS_NOR2X2 U14320 ( .A(n6175), .B(n6269), .Z(n6626) );
  HS65_LS_NOR2X2 U14321 ( .A(n3147), .B(n3173), .Z(n3762) );
  HS65_LS_NOR2X2 U14322 ( .A(n1312), .B(n1208), .Z(n1226) );
  HS65_LS_NOR2X2 U14323 ( .A(n6481), .B(n6529), .Z(n6512) );
  HS65_LS_NOR2X2 U14324 ( .A(n6595), .B(n6583), .Z(n6566) );
  HS65_LS_NOR2X2 U14325 ( .A(n5002), .B(n4990), .Z(n4973) );
  HS65_LS_NOR2X2 U14326 ( .A(n4888), .B(n4936), .Z(n4919) );
  HS65_LS_NOR2X2 U14327 ( .A(n4874), .B(n4861), .Z(n4843) );
  HS65_LS_NOR2X2 U14328 ( .A(n6467), .B(n6454), .Z(n6436) );
  HS65_LS_NOR2X2 U14329 ( .A(n7953), .B(n7954), .Z(n8586) );
  HS65_LS_NAND2X2 U14330 ( .A(n6170), .B(n6087), .Z(n6679) );
  HS65_LS_NAND2X2 U14331 ( .A(n4577), .B(n4494), .Z(n5086) );
  HS65_LS_NOR2AX3 U14332 ( .A(n4616), .B(n4509), .Z(n5415) );
  HS65_LS_NOR2AX3 U14333 ( .A(n4591), .B(n4463), .Z(n5300) );
  HS65_LS_NOR2AX3 U14334 ( .A(n6209), .B(n6102), .Z(n7007) );
  HS65_LS_NOR2AX3 U14335 ( .A(n4531), .B(n4862), .Z(n5184) );
  HS65_LS_NOR2AX3 U14336 ( .A(n6184), .B(n6056), .Z(n6892) );
  HS65_LS_NOR2AX3 U14337 ( .A(n6124), .B(n6455), .Z(n6776) );
  HS65_LS_NOR2X2 U14338 ( .A(n8004), .B(n7871), .Z(n8300) );
  HS65_LS_NOR2X2 U14339 ( .A(n2064), .B(n1960), .Z(n1978) );
  HS65_LS_NOR2X2 U14340 ( .A(n3625), .B(n3585), .Z(n3598) );
  HS65_LS_NOR2X2 U14341 ( .A(n4669), .B(n4721), .Z(n4703) );
  HS65_LS_NOR2X2 U14342 ( .A(n6262), .B(n6314), .Z(n6296) );
  HS65_LS_NOR2X2 U14343 ( .A(n3728), .B(n3353), .Z(n3312) );
  HS65_LS_NOR2X2 U14344 ( .A(n1154), .B(n1201), .Z(n1241) );
  HS65_LS_NOR2X2 U14345 ( .A(n1906), .B(n1953), .Z(n1993) );
  HS65_LS_NOR2X2 U14346 ( .A(n1530), .B(n1577), .Z(n1617) );
  HS65_LS_NOR2X2 U14347 ( .A(n2282), .B(n2329), .Z(n2369) );
  HS65_LS_NAND2X2 U14348 ( .A(n8164), .B(n7846), .Z(n8400) );
  HS65_LS_NAND2X2 U14349 ( .A(n8196), .B(n7885), .Z(n8460) );
  HS65_LS_NOR2X2 U14350 ( .A(n3282), .B(n3065), .Z(n3641) );
  HS65_LS_NAND2X2 U14351 ( .A(n7818), .B(n7978), .Z(n7815) );
  HS65_LS_NAND2X2 U14352 ( .A(n7917), .B(n7991), .Z(n7915) );
  HS65_LS_NAND2X2 U14353 ( .A(n8542), .B(n7961), .Z(n8365) );
  HS65_LS_NOR2X2 U14354 ( .A(n7978), .B(n7686), .Z(n8408) );
  HS65_LS_NOR2X2 U14355 ( .A(n7991), .B(n7724), .Z(n8468) );
  HS65_LS_NOR2X2 U14356 ( .A(n4495), .B(n5524), .Z(n5056) );
  HS65_LS_NOR2X2 U14357 ( .A(n6088), .B(n7116), .Z(n6649) );
  HS65_LS_NOR2X2 U14358 ( .A(n1548), .B(n1775), .Z(n1722) );
  HS65_LS_NOR2X2 U14359 ( .A(n2300), .B(n2527), .Z(n2474) );
  HS65_LS_NOR2X2 U14360 ( .A(n6064), .B(n6337), .Z(n6884) );
  HS65_LS_NOR2X2 U14361 ( .A(n4471), .B(n4744), .Z(n5292) );
  HS65_LS_NOR2X2 U14362 ( .A(n4517), .B(n4783), .Z(n5407) );
  HS65_LS_NOR2X2 U14363 ( .A(n6110), .B(n6376), .Z(n6999) );
  HS65_LS_NOR2X2 U14364 ( .A(n5508), .B(n4637), .Z(n5175) );
  HS65_LS_NOR2X2 U14365 ( .A(n7100), .B(n6230), .Z(n6767) );
  HS65_LS_NOR2X2 U14366 ( .A(n3280), .B(n3063), .Z(n3593) );
  HS65_LS_NOR2X2 U14367 ( .A(n6056), .B(n6058), .Z(n6864) );
  HS65_LS_NOR2X2 U14368 ( .A(n4463), .B(n4465), .Z(n5272) );
  HS65_LS_NOR2X2 U14369 ( .A(n4509), .B(n4511), .Z(n5387) );
  HS65_LS_NOR2X2 U14370 ( .A(n6102), .B(n6104), .Z(n6979) );
  HS65_LS_NOR2X2 U14371 ( .A(n4862), .B(n4636), .Z(n5155) );
  HS65_LS_NOR2X2 U14372 ( .A(n6455), .B(n6229), .Z(n6747) );
  HS65_LS_NOR2X2 U14373 ( .A(n3007), .B(n3983), .Z(n3418) );
  HS65_LS_NOR2X2 U14374 ( .A(n7846), .B(n7638), .Z(n7808) );
  HS65_LS_NOR2X2 U14375 ( .A(n7885), .B(n7666), .Z(n7908) );
  HS65_LS_NOR2X2 U14376 ( .A(n3985), .B(n3391), .Z(n3385) );
  HS65_LS_NOR2X2 U14377 ( .A(n7857), .B(n7869), .Z(n8117) );
  HS65_LS_NOR2X2 U14378 ( .A(n1172), .B(n1399), .Z(n1346) );
  HS65_LS_NOR2X2 U14379 ( .A(n8051), .B(n8045), .Z(n8550) );
  HS65_LS_NOR2X2 U14380 ( .A(n8045), .B(n8361), .Z(n8615) );
  HS65_LS_NOR2X2 U14381 ( .A(n4503), .B(n4613), .Z(n5434) );
  HS65_LS_NOR2X2 U14382 ( .A(n4457), .B(n4601), .Z(n5319) );
  HS65_LS_NOR2X2 U14383 ( .A(n4835), .B(n4543), .Z(n5203) );
  HS65_LS_NOR2X2 U14384 ( .A(n6096), .B(n6206), .Z(n7026) );
  HS65_LS_NOR2X2 U14385 ( .A(n6050), .B(n6194), .Z(n6911) );
  HS65_LS_NOR2X2 U14386 ( .A(n6428), .B(n6136), .Z(n6795) );
  HS65_LS_NOR2X2 U14387 ( .A(n1505), .B(n1571), .Z(n1726) );
  HS65_LS_NOR2X2 U14388 ( .A(n2257), .B(n2323), .Z(n2478) );
  HS65_LS_NOR2X2 U14389 ( .A(n8671), .B(n8030), .Z(n8113) );
  HS65_LS_NOR2X2 U14390 ( .A(n1924), .B(n2151), .Z(n2098) );
  HS65_LS_NOR2X2 U14391 ( .A(n3262), .B(n3057), .Z(n3563) );
  HS65_LS_NOR2X2 U14392 ( .A(n7210), .B(n7204), .Z(n6873) );
  HS65_LS_NOR2X2 U14393 ( .A(n5618), .B(n5612), .Z(n5281) );
  HS65_LS_NOR2X2 U14394 ( .A(n5645), .B(n5639), .Z(n5396) );
  HS65_LS_NOR2X2 U14395 ( .A(n7237), .B(n7231), .Z(n6988) );
  HS65_LS_NOR2X2 U14396 ( .A(n5591), .B(n5588), .Z(n5164) );
  HS65_LS_NOR2X2 U14397 ( .A(n7183), .B(n7180), .Z(n6756) );
  HS65_LS_NAND2X2 U14398 ( .A(n3585), .B(n2925), .Z(n3268) );
  HS65_LS_NOR2X2 U14399 ( .A(n1128), .B(n1376), .Z(n1285) );
  HS65_LS_NOR2X2 U14400 ( .A(n1880), .B(n2128), .Z(n2037) );
  HS65_LS_NOR2X2 U14401 ( .A(n2256), .B(n2504), .Z(n2413) );
  HS65_LS_NOR2X2 U14402 ( .A(n1504), .B(n1752), .Z(n1661) );
  HS65_LS_NOR2X2 U14403 ( .A(n4516), .B(n5565), .Z(n5410) );
  HS65_LS_NOR2X2 U14404 ( .A(n4470), .B(n5544), .Z(n5295) );
  HS65_LS_NOR2X2 U14405 ( .A(n4535), .B(n5589), .Z(n5178) );
  HS65_LS_NOR2X2 U14406 ( .A(n6109), .B(n7157), .Z(n7002) );
  HS65_LS_NOR2X2 U14407 ( .A(n6063), .B(n7136), .Z(n6887) );
  HS65_LS_NOR2X2 U14408 ( .A(n6128), .B(n7181), .Z(n6770) );
  HS65_LS_NAND2X2 U14409 ( .A(n8182), .B(n8181), .Z(n7748) );
  HS65_LS_NAND2X2 U14410 ( .A(n8150), .B(n8149), .Z(n7710) );
  HS65_LS_NAND2X2 U14411 ( .A(n6153), .B(n6313), .Z(n6172) );
  HS65_LS_NAND2X2 U14412 ( .A(n4560), .B(n4720), .Z(n4579) );
  HS65_LS_NAND2X2 U14413 ( .A(n6058), .B(n6528), .Z(n6356) );
  HS65_LS_NAND2X2 U14414 ( .A(n4465), .B(n4935), .Z(n4763) );
  HS65_LS_NAND2X2 U14415 ( .A(n4511), .B(n4989), .Z(n4802) );
  HS65_LS_NAND2X2 U14416 ( .A(n6104), .B(n6582), .Z(n6395) );
  HS65_LS_NAND2X2 U14417 ( .A(n6229), .B(n6452), .Z(n6249) );
  HS65_LS_NAND2X2 U14418 ( .A(n4636), .B(n4859), .Z(n4656) );
  HS65_LS_NAND2X2 U14419 ( .A(n3053), .B(n4103), .Z(n3608) );
  HS65_LS_NOR2X2 U14420 ( .A(n1129), .B(n1195), .Z(n1350) );
  HS65_LS_NOR2X2 U14421 ( .A(n1881), .B(n1947), .Z(n2102) );
  HS65_LS_NOR2X2 U14422 ( .A(n1404), .B(n1243), .Z(n1237) );
  HS65_LS_NOR2X2 U14423 ( .A(n2156), .B(n1995), .Z(n1989) );
  HS65_LS_NOR2X2 U14424 ( .A(n2532), .B(n2371), .Z(n2365) );
  HS65_LS_NOR2X2 U14425 ( .A(n1780), .B(n1619), .Z(n1613) );
  HS65_LS_NOR2X2 U14426 ( .A(n8003), .B(n8119), .Z(n8236) );
  HS65_LS_NOR2X2 U14427 ( .A(n4488), .B(n5517), .Z(n5108) );
  HS65_LS_NOR2X2 U14428 ( .A(n6081), .B(n7109), .Z(n6701) );
  HS65_LS_NOR2X2 U14429 ( .A(n7959), .B(n7779), .Z(n8582) );
  HS65_LS_NOR2X2 U14430 ( .A(n7857), .B(n7762), .Z(n8278) );
  HS65_LS_NOR2X2 U14431 ( .A(n4562), .B(n5524), .Z(n5073) );
  HS65_LS_NOR2X2 U14432 ( .A(n6155), .B(n7116), .Z(n6666) );
  HS65_LS_NOR2X2 U14433 ( .A(n6315), .B(n6153), .Z(n6627) );
  HS65_LS_NOR2X2 U14434 ( .A(n4722), .B(n4560), .Z(n5034) );
  HS65_LS_NOR2X2 U14435 ( .A(n7646), .B(n7638), .Z(n8723) );
  HS65_LS_NOR2X2 U14436 ( .A(n7674), .B(n7666), .Z(n8811) );
  HS65_LS_NOR2X2 U14437 ( .A(n2971), .B(n2965), .Z(n3479) );
  HS65_LS_NOR2X2 U14438 ( .A(n3964), .B(n3329), .Z(n3323) );
  HS65_LS_NOR2X2 U14439 ( .A(n3262), .B(n2927), .Z(n3646) );
  HS65_LS_NOR2X2 U14440 ( .A(n3905), .B(n3536), .Z(n3531) );
  HS65_LS_NOR2X2 U14441 ( .A(n7632), .B(n7847), .Z(n8410) );
  HS65_LS_NOR2X2 U14442 ( .A(n7660), .B(n7886), .Z(n8470) );
  HS65_LS_NOR2X2 U14443 ( .A(n7870), .B(n7871), .Z(n8282) );
  HS65_LS_NOR2X2 U14444 ( .A(n1780), .B(n1530), .Z(n1689) );
  HS65_LS_NOR2X2 U14445 ( .A(n2532), .B(n2282), .Z(n2441) );
  HS65_LS_NOR2X2 U14446 ( .A(n6051), .B(n7204), .Z(n6952) );
  HS65_LS_NOR2X2 U14447 ( .A(n6097), .B(n7231), .Z(n7067) );
  HS65_LS_NOR2X2 U14448 ( .A(n4504), .B(n5639), .Z(n5475) );
  HS65_LS_NOR2X2 U14449 ( .A(n4458), .B(n5612), .Z(n5360) );
  HS65_LS_NOR2X2 U14450 ( .A(n4820), .B(n5588), .Z(n5245) );
  HS65_LS_NOR2X2 U14451 ( .A(n6413), .B(n7180), .Z(n6837) );
  HS65_LS_NOR2X2 U14452 ( .A(n3101), .B(n2961), .Z(n3446) );
  HS65_LS_NOR2X2 U14453 ( .A(n1511), .B(n1752), .Z(n1748) );
  HS65_LS_NOR2X2 U14454 ( .A(n2263), .B(n2504), .Z(n2500) );
  HS65_LS_NOR2X2 U14455 ( .A(n1135), .B(n1376), .Z(n1372) );
  HS65_LS_NOR2X2 U14456 ( .A(n1887), .B(n2128), .Z(n2124) );
  HS65_LS_NOR2X2 U14457 ( .A(n4559), .B(n4487), .Z(n5112) );
  HS65_LS_NOR2X2 U14458 ( .A(n6152), .B(n6080), .Z(n6705) );
  HS65_LS_NOR2X2 U14459 ( .A(n7960), .B(n8051), .Z(n8605) );
  HS65_LS_NAND2X2 U14460 ( .A(n2943), .B(n2874), .Z(n2963) );
  HS65_LS_NOR2X2 U14461 ( .A(n1404), .B(n1154), .Z(n1313) );
  HS65_LS_NOR2X2 U14462 ( .A(n2156), .B(n1906), .Z(n2065) );
  HS65_LS_NOR2X2 U14463 ( .A(n2257), .B(n2328), .Z(n2410) );
  HS65_LS_NOR2X2 U14464 ( .A(n1505), .B(n1576), .Z(n1658) );
  HS65_LS_NAND2X2 U14465 ( .A(n2255), .B(n2250), .Z(n2345) );
  HS65_LS_NAND2X2 U14466 ( .A(n1127), .B(n1122), .Z(n1217) );
  HS65_LS_NAND2X2 U14467 ( .A(n1879), .B(n1874), .Z(n1969) );
  HS65_LS_NAND2X2 U14468 ( .A(n1503), .B(n1498), .Z(n1593) );
  HS65_LS_NOR2X2 U14469 ( .A(n7817), .B(n7635), .Z(n7802) );
  HS65_LS_NOR2X2 U14470 ( .A(n7880), .B(n7663), .Z(n7902) );
  HS65_LS_NOR2X2 U14471 ( .A(n2849), .B(n3203), .Z(n3883) );
  HS65_LS_NOR2AX3 U14472 ( .A(n7709), .B(n7687), .Z(n8711) );
  HS65_LS_NOR2AX3 U14473 ( .A(n7747), .B(n7725), .Z(n8799) );
  HS65_LS_NOR2X2 U14474 ( .A(n7084), .B(n7109), .Z(n6714) );
  HS65_LS_NOR2X2 U14475 ( .A(n5492), .B(n5517), .Z(n5121) );
  HS65_LS_NOR2X2 U14476 ( .A(n4799), .B(n5009), .Z(n4988) );
  HS65_LS_NOR2X2 U14477 ( .A(n4760), .B(n4895), .Z(n4934) );
  HS65_LS_NOR2X2 U14478 ( .A(n6392), .B(n6602), .Z(n6581) );
  HS65_LS_NOR2X2 U14479 ( .A(n4576), .B(n4677), .Z(n4718) );
  HS65_LS_NOR2X2 U14480 ( .A(n6353), .B(n6488), .Z(n6527) );
  HS65_LS_NOR2X2 U14481 ( .A(n6169), .B(n6270), .Z(n6311) );
  HS65_LS_NOR2X2 U14482 ( .A(n4653), .B(n4881), .Z(n4858) );
  HS65_LS_NOR2X2 U14483 ( .A(n6246), .B(n6474), .Z(n6451) );
  HS65_LS_NOR2X2 U14484 ( .A(n7959), .B(n7952), .Z(n8359) );
  HS65_LS_NOR2X2 U14485 ( .A(n1129), .B(n1200), .Z(n1282) );
  HS65_LS_NOR2X2 U14486 ( .A(n1881), .B(n1952), .Z(n2034) );
  HS65_LS_NOR2X2 U14487 ( .A(n3942), .B(n2873), .Z(n3487) );
  HS65_LS_NOR2X2 U14488 ( .A(n8030), .B(n8009), .Z(n8104) );
  HS65_LS_NOR2X2 U14489 ( .A(n3174), .B(n3147), .Z(n3720) );
  HS65_LS_NOR2X2 U14490 ( .A(n2849), .B(n3208), .Z(n3799) );
  HS65_LS_NAND2X2 U14491 ( .A(n7660), .B(n8472), .Z(n8194) );
  HS65_LS_NAND2X2 U14492 ( .A(n7632), .B(n8412), .Z(n8162) );
  HS65_LS_NOR2X2 U14493 ( .A(n8335), .B(n7955), .Z(n8366) );
  HS65_LS_NAND2X2 U14494 ( .A(n2895), .B(n2986), .Z(n3165) );
  HS65_LS_NOR2X2 U14495 ( .A(n6155), .B(n6262), .Z(n6676) );
  HS65_LS_NOR2X2 U14496 ( .A(n4562), .B(n4669), .Z(n5083) );
  HS65_LS_NOR2X2 U14497 ( .A(n8881), .B(n8069), .Z(n8355) );
  HS65_LS_NOR2X2 U14498 ( .A(n6358), .B(n6065), .Z(n6913) );
  HS65_LS_NOR2X2 U14499 ( .A(n4765), .B(n4472), .Z(n5321) );
  HS65_LS_NOR2X2 U14500 ( .A(n4804), .B(n4518), .Z(n5436) );
  HS65_LS_NOR2X2 U14501 ( .A(n6397), .B(n6111), .Z(n7028) );
  HS65_LS_NOR2X2 U14502 ( .A(n4658), .B(n4533), .Z(n5205) );
  HS65_LS_NOR2X2 U14503 ( .A(n6251), .B(n6126), .Z(n6797) );
  HS65_LS_NAND2X2 U14504 ( .A(n4800), .B(n4618), .Z(n5439) );
  HS65_LS_NAND2X2 U14505 ( .A(n4761), .B(n4593), .Z(n5324) );
  HS65_LS_NAND2X2 U14506 ( .A(n4654), .B(n4534), .Z(n5208) );
  HS65_LS_NAND2X2 U14507 ( .A(n6393), .B(n6211), .Z(n7031) );
  HS65_LS_NAND2X2 U14508 ( .A(n6354), .B(n6186), .Z(n6916) );
  HS65_LS_NAND2X2 U14509 ( .A(n6247), .B(n6127), .Z(n6800) );
  HS65_LS_NAND2X2 U14510 ( .A(n3044), .B(n3043), .Z(n3050) );
  HS65_LS_NOR2X2 U14511 ( .A(n3003), .B(n3209), .Z(n3389) );
  HS65_LS_NOR2X2 U14512 ( .A(n2873), .B(n2966), .Z(n3098) );
  HS65_LS_NOR2X2 U14513 ( .A(n3985), .B(n3003), .Z(n3846) );
  HS65_LS_NOR2X2 U14514 ( .A(n4989), .B(n4503), .Z(n5478) );
  HS65_LS_NOR2X2 U14515 ( .A(n4935), .B(n4457), .Z(n5363) );
  HS65_LS_NOR2X2 U14516 ( .A(n6582), .B(n6096), .Z(n7070) );
  HS65_LS_NOR2X2 U14517 ( .A(n6528), .B(n6050), .Z(n6955) );
  HS65_LS_NOR2X2 U14518 ( .A(n4859), .B(n4835), .Z(n5248) );
  HS65_LS_NOR2X2 U14519 ( .A(n6452), .B(n6428), .Z(n6840) );
  HS65_LS_NOR2X2 U14520 ( .A(n7885), .B(n7663), .Z(n8835) );
  HS65_LS_NOR2X2 U14521 ( .A(n7846), .B(n7635), .Z(n8747) );
  HS65_LS_NOR2X2 U14522 ( .A(n8030), .B(n7999), .Z(n8232) );
  HS65_LS_NOR2X2 U14523 ( .A(n7846), .B(n8149), .Z(n8708) );
  HS65_LS_NOR2X2 U14524 ( .A(n7885), .B(n8181), .Z(n8796) );
  HS65_LS_NAND2X2 U14525 ( .A(n2961), .B(n3942), .Z(n3467) );
  HS65_LS_NOR2X2 U14526 ( .A(n2986), .B(n3174), .Z(n3763) );
  HS65_LS_NAND2X2 U14527 ( .A(n1572), .B(n1780), .Z(n1732) );
  HS65_LS_NAND2X2 U14528 ( .A(n2324), .B(n2532), .Z(n2484) );
  HS65_LS_NOR2X2 U14529 ( .A(n4785), .B(n5565), .Z(n5426) );
  HS65_LS_NOR2X2 U14530 ( .A(n4746), .B(n5544), .Z(n5311) );
  HS65_LS_NOR2X2 U14531 ( .A(n6378), .B(n7157), .Z(n7018) );
  HS65_LS_NOR2X2 U14532 ( .A(n4639), .B(n5589), .Z(n5195) );
  HS65_LS_NOR2X2 U14533 ( .A(n6232), .B(n7181), .Z(n6787) );
  HS65_LS_NOR2X2 U14534 ( .A(n6339), .B(n7136), .Z(n6903) );
  HS65_LS_AOI212X2 U14535 ( .A(n152), .B(n3608), .C(n156), .D(n176), .E(n4121), 
        .Z(n4118) );
  HS65_LS_CBI4I1X3 U14536 ( .A(n3045), .B(n2928), .C(n3053), .D(n3554), .Z(
        n4121) );
  HS65_LS_NAND2X2 U14537 ( .A(n3208), .B(n2855), .Z(n3376) );
  HS65_LS_NOR2X2 U14538 ( .A(n5526), .B(n5523), .Z(n5042) );
  HS65_LS_NOR2X2 U14539 ( .A(n7118), .B(n7115), .Z(n6635) );
  HS65_LS_NOR2X2 U14540 ( .A(n8060), .B(n7963), .Z(n8621) );
  HS65_LS_NOR4ABX2 U14541 ( .A(n3998), .B(n3999), .C(n4000), .D(n4001), .Z(
        n3925) );
  HS65_LS_OAI222X2 U14542 ( .A(n4002), .B(n3599), .C(n3065), .D(n2924), .E(
        n3045), .F(n3280), .Z(n4001) );
  HS65_LS_OAI212X3 U14543 ( .A(n3586), .B(n3067), .C(n2925), .D(n3263), .E(
        n4003), .Z(n4000) );
  HS65_LS_NOR3AX2 U14544 ( .A(n3254), .B(n3567), .C(n3041), .Z(n3998) );
  HS65_LS_NAND2X2 U14545 ( .A(n1948), .B(n2156), .Z(n2108) );
  HS65_LS_NAND2X2 U14546 ( .A(n1196), .B(n1404), .Z(n1356) );
  HS65_LS_NOR2X2 U14547 ( .A(n8149), .B(n7697), .Z(n8763) );
  HS65_LS_NOR2X2 U14548 ( .A(n8181), .B(n7735), .Z(n8851) );
  HS65_LS_NOR4ABX2 U14549 ( .A(n1800), .B(n1801), .C(n1802), .D(n1803), .Z(
        n1765) );
  HS65_LS_OAI222X2 U14550 ( .A(n1776), .B(n1529), .C(n1775), .D(n1531), .E(
        n1686), .F(n1548), .Z(n1803) );
  HS65_LS_NOR3X1 U14551 ( .A(n1666), .B(n1551), .C(n1620), .Z(n1800) );
  HS65_LS_OAI212X3 U14552 ( .A(n1753), .B(n1497), .C(n1532), .D(n1619), .E(
        n1804), .Z(n1802) );
  HS65_LS_NOR4ABX2 U14553 ( .A(n2552), .B(n2553), .C(n2554), .D(n2555), .Z(
        n2517) );
  HS65_LS_OAI222X2 U14554 ( .A(n2528), .B(n2281), .C(n2527), .D(n2283), .E(
        n2438), .F(n2300), .Z(n2555) );
  HS65_LS_NOR3X1 U14555 ( .A(n2418), .B(n2303), .C(n2372), .Z(n2552) );
  HS65_LS_OAI212X3 U14556 ( .A(n2505), .B(n2249), .C(n2284), .D(n2371), .E(
        n2556), .Z(n2554) );
  HS65_LS_NOR4ABX2 U14557 ( .A(n1424), .B(n1425), .C(n1426), .D(n1427), .Z(
        n1389) );
  HS65_LS_OAI222X2 U14558 ( .A(n1400), .B(n1153), .C(n1399), .D(n1155), .E(
        n1310), .F(n1172), .Z(n1427) );
  HS65_LS_NOR3X1 U14559 ( .A(n1290), .B(n1175), .C(n1244), .Z(n1424) );
  HS65_LS_OAI212X3 U14560 ( .A(n1377), .B(n1121), .C(n1156), .D(n1243), .E(
        n1428), .Z(n1426) );
  HS65_LS_NOR4ABX2 U14561 ( .A(n2176), .B(n2177), .C(n2178), .D(n2179), .Z(
        n2141) );
  HS65_LS_OAI222X2 U14562 ( .A(n2152), .B(n1905), .C(n2151), .D(n1907), .E(
        n2062), .F(n1924), .Z(n2179) );
  HS65_LS_NOR3X1 U14563 ( .A(n2042), .B(n1927), .C(n1996), .Z(n2176) );
  HS65_LS_OAI212X3 U14564 ( .A(n2129), .B(n1873), .C(n1908), .D(n1995), .E(
        n2180), .Z(n2178) );
  HS65_LS_NOR2X2 U14565 ( .A(n3391), .B(n3215), .Z(n3375) );
  HS65_LS_NOR2X2 U14566 ( .A(n3329), .B(n3163), .Z(n3690) );
  HS65_LS_NOR2X2 U14567 ( .A(n7109), .B(n7118), .Z(n6688) );
  HS65_LS_NOR2X2 U14568 ( .A(n5517), .B(n5526), .Z(n5095) );
  HS65_LS_NOR2X2 U14569 ( .A(n4504), .B(n4800), .Z(n5411) );
  HS65_LS_NOR2X2 U14570 ( .A(n4458), .B(n4761), .Z(n5296) );
  HS65_LS_NOR2X2 U14571 ( .A(n6097), .B(n6393), .Z(n7003) );
  HS65_LS_NOR2X2 U14572 ( .A(n4820), .B(n4654), .Z(n5179) );
  HS65_LS_NOR2X2 U14573 ( .A(n6051), .B(n6354), .Z(n6888) );
  HS65_LS_NOR2X2 U14574 ( .A(n6413), .B(n6247), .Z(n6771) );
  HS65_LS_NOR2X2 U14575 ( .A(n1619), .B(n1572), .Z(n1666) );
  HS65_LS_NOR2X2 U14576 ( .A(n2371), .B(n2324), .Z(n2418) );
  HS65_LS_NOR2X2 U14577 ( .A(n3895), .B(n2849), .Z(n3407) );
  HS65_LS_NAND2X2 U14578 ( .A(n1130), .B(n1155), .Z(n1198) );
  HS65_LS_NAND2X2 U14579 ( .A(n1882), .B(n1907), .Z(n1950) );
  HS65_LS_NAND2X2 U14580 ( .A(n2258), .B(n2283), .Z(n2326) );
  HS65_LS_NAND2X2 U14581 ( .A(n1506), .B(n1531), .Z(n1574) );
  HS65_LS_NOR2X2 U14582 ( .A(n1995), .B(n1948), .Z(n2042) );
  HS65_LS_NOR2X2 U14583 ( .A(n1243), .B(n1196), .Z(n1290) );
  HS65_LS_NOR2X2 U14584 ( .A(n4680), .B(n5523), .Z(n5109) );
  HS65_LS_NOR2X2 U14585 ( .A(n6273), .B(n7115), .Z(n6702) );
  HS65_LS_NOR2X2 U14586 ( .A(n3263), .B(n3290), .Z(n3245) );
  HS65_LS_NOR2X2 U14587 ( .A(n3391), .B(n3204), .Z(n3807) );
  HS65_LS_NOR2X2 U14588 ( .A(n3625), .B(n3044), .Z(n3040) );
  HS65_LS_NOR4ABX2 U14589 ( .A(n2295), .B(n2296), .C(n2297), .D(n2298), .Z(
        n2275) );
  HS65_LS_OAI212X3 U14590 ( .A(n2258), .B(n2299), .C(n2300), .D(n2301), .E(
        n2302), .Z(n2298) );
  HS65_LS_NOR4ABX2 U14591 ( .A(n2307), .B(n2308), .C(n2309), .D(n2310), .Z(
        n2296) );
  HS65_LS_NOR3AX2 U14592 ( .A(n2311), .B(n2312), .C(n2313), .Z(n2295) );
  HS65_LS_NOR4ABX2 U14593 ( .A(n1543), .B(n1544), .C(n1545), .D(n1546), .Z(
        n1523) );
  HS65_LS_OAI212X3 U14594 ( .A(n1506), .B(n1547), .C(n1548), .D(n1549), .E(
        n1550), .Z(n1546) );
  HS65_LS_NOR4ABX2 U14595 ( .A(n1555), .B(n1556), .C(n1557), .D(n1558), .Z(
        n1544) );
  HS65_LS_NOR3AX2 U14596 ( .A(n1559), .B(n1560), .C(n1561), .Z(n1543) );
  HS65_LS_NOR4ABX2 U14597 ( .A(n1167), .B(n1168), .C(n1169), .D(n1170), .Z(
        n1147) );
  HS65_LS_OAI212X3 U14598 ( .A(n1130), .B(n1171), .C(n1172), .D(n1173), .E(
        n1174), .Z(n1170) );
  HS65_LS_NOR3AX2 U14599 ( .A(n1183), .B(n1184), .C(n1185), .Z(n1167) );
  HS65_LS_NOR4ABX2 U14600 ( .A(n1179), .B(n1180), .C(n1181), .D(n1182), .Z(
        n1168) );
  HS65_LS_NOR4ABX2 U14601 ( .A(n1919), .B(n1920), .C(n1921), .D(n1922), .Z(
        n1899) );
  HS65_LS_OAI212X3 U14602 ( .A(n1882), .B(n1923), .C(n1924), .D(n1925), .E(
        n1926), .Z(n1922) );
  HS65_LS_NOR3AX2 U14603 ( .A(n1935), .B(n1936), .C(n1937), .Z(n1919) );
  HS65_LS_NOR4ABX2 U14604 ( .A(n1931), .B(n1932), .C(n1933), .D(n1934), .Z(
        n1920) );
  HS65_LS_NOR2X2 U14605 ( .A(n2923), .B(n3044), .Z(n3037) );
  HS65_LS_NOR2X2 U14606 ( .A(n8069), .B(n8041), .Z(n8619) );
  HS65_LS_NOR2X2 U14607 ( .A(n3964), .B(n2985), .Z(n3729) );
  HS65_LS_NAND2X2 U14608 ( .A(n8041), .B(n8881), .Z(n8553) );
  HS65_LS_NOR2X2 U14609 ( .A(n4576), .B(n4719), .Z(n5081) );
  HS65_LS_NOR2X2 U14610 ( .A(n6169), .B(n6312), .Z(n6674) );
  HS65_LS_NOR2X2 U14611 ( .A(n2873), .B(n2946), .Z(n2954) );
  HS65_LS_NAND2X2 U14612 ( .A(n3042), .B(n2924), .Z(n3055) );
  HS65_LS_NOR2X2 U14613 ( .A(n6358), .B(n6488), .Z(n6906) );
  HS65_LS_NOR2X2 U14614 ( .A(n6174), .B(n6270), .Z(n6669) );
  HS65_LS_NOR2X2 U14615 ( .A(n4581), .B(n4677), .Z(n5076) );
  HS65_LS_NOR2X2 U14616 ( .A(n4804), .B(n5009), .Z(n5429) );
  HS65_LS_NOR2X2 U14617 ( .A(n6397), .B(n6602), .Z(n7021) );
  HS65_LS_NOR2X2 U14618 ( .A(n4765), .B(n4895), .Z(n5314) );
  HS65_LS_NOR2X2 U14619 ( .A(n4658), .B(n4881), .Z(n5198) );
  HS65_LS_NOR2X2 U14620 ( .A(n6251), .B(n6474), .Z(n6790) );
  HS65_LS_NOR2X2 U14621 ( .A(n8332), .B(n8639), .Z(n8609) );
  HS65_LS_NAND2X2 U14622 ( .A(n3163), .B(n3964), .Z(n3710) );
  HS65_LS_NOR2X2 U14623 ( .A(n7191), .B(n7210), .Z(n6925) );
  HS65_LS_NOR2X2 U14624 ( .A(n5599), .B(n5618), .Z(n5333) );
  HS65_LS_NOR2X2 U14625 ( .A(n5626), .B(n5645), .Z(n5448) );
  HS65_LS_NOR2X2 U14626 ( .A(n7218), .B(n7237), .Z(n7040) );
  HS65_LS_NOR2X2 U14627 ( .A(n7174), .B(n7183), .Z(n6809) );
  HS65_LS_NOR2X2 U14628 ( .A(n5582), .B(n5591), .Z(n5217) );
  HS65_LS_NOR2X2 U14629 ( .A(n7847), .B(n8164), .Z(n8729) );
  HS65_LS_NOR2X2 U14630 ( .A(n7886), .B(n8196), .Z(n8817) );
  HS65_LS_NOR2X2 U14631 ( .A(n2877), .B(n3940), .Z(n3130) );
  HS65_LS_NOR2X2 U14632 ( .A(n2966), .B(n3470), .Z(n3503) );
  HS65_LS_NOR2X2 U14633 ( .A(n3065), .B(n3052), .Z(n3555) );
  HS65_LS_NAND2X2 U14634 ( .A(n7999), .B(n8671), .Z(n8249) );
  HS65_LS_NAND2X2 U14635 ( .A(n4618), .B(n5009), .Z(n4523) );
  HS65_LS_NAND2X2 U14636 ( .A(n6211), .B(n6602), .Z(n6116) );
  HS65_LS_NAND2X2 U14637 ( .A(n6186), .B(n6488), .Z(n6070) );
  HS65_LS_NAND2X2 U14638 ( .A(n4593), .B(n4895), .Z(n4477) );
  HS65_LS_NAND2X2 U14639 ( .A(n6127), .B(n6474), .Z(n7097) );
  HS65_LS_NAND2X2 U14640 ( .A(n4494), .B(n4677), .Z(n5489) );
  HS65_LS_NAND2X2 U14641 ( .A(n6087), .B(n6270), .Z(n7081) );
  HS65_LS_NAND2X2 U14642 ( .A(n4534), .B(n4881), .Z(n5505) );
  HS65_LS_NOR2X2 U14643 ( .A(n7952), .B(n8556), .Z(n8585) );
  HS65_LS_NOR2X2 U14644 ( .A(n7869), .B(n8252), .Z(n8281) );
  HS65_LS_NOR2X2 U14645 ( .A(n4002), .B(n2927), .Z(n3294) );
  HS65_LS_NOR2X2 U14646 ( .A(n8018), .B(n7861), .Z(n8230) );
  HS65_LS_CBI4I1X3 U14647 ( .A(n1506), .B(n1534), .C(n1584), .D(n1664), .Z(
        n1818) );
  HS65_LS_CBI4I1X3 U14648 ( .A(n2258), .B(n2286), .C(n2336), .D(n2416), .Z(
        n2570) );
  HS65_LS_CBI4I1X3 U14649 ( .A(n3290), .B(n3044), .C(n3063), .D(n3611), .Z(
        n3610) );
  HS65_LS_CBI4I1X3 U14650 ( .A(n3127), .B(n2946), .C(n3470), .D(n3471), .Z(
        n3469) );
  HS65_LS_NOR2X2 U14651 ( .A(n2256), .B(n2336), .Z(n2400) );
  HS65_LS_NOR2X2 U14652 ( .A(n1504), .B(n1584), .Z(n1648) );
  HS65_LS_CBI4I1X3 U14653 ( .A(n1130), .B(n1158), .C(n1208), .D(n1288), .Z(
        n1442) );
  HS65_LS_NOR2X2 U14654 ( .A(n3778), .B(n2894), .Z(n3345) );
  HS65_LS_NOR2X2 U14655 ( .A(n3538), .B(n3100), .Z(n3118) );
  HS65_LS_NOR2X2 U14656 ( .A(n2985), .B(n3148), .Z(n3156) );
  HS65_LS_NOR2X2 U14657 ( .A(n1128), .B(n1208), .Z(n1272) );
  HS65_LS_NOR2X2 U14658 ( .A(n2257), .B(n2286), .Z(n2454) );
  HS65_LS_NOR2X2 U14659 ( .A(n1505), .B(n1534), .Z(n1702) );
  HS65_LS_CBI4I1X3 U14660 ( .A(n1882), .B(n1910), .C(n1960), .D(n2040), .Z(
        n2194) );
  HS65_LS_NAND2X2 U14661 ( .A(n3625), .B(n2924), .Z(n3552) );
  HS65_LS_CBI4I1X3 U14662 ( .A(n2895), .B(n2989), .C(n3353), .D(n3688), .Z(
        n4246) );
  HS65_LS_NOR2X2 U14663 ( .A(n2282), .B(n2528), .Z(n2442) );
  HS65_LS_NOR2X2 U14664 ( .A(n1530), .B(n1776), .Z(n1690) );
  HS65_LS_NAND2X2 U14665 ( .A(n3895), .B(n2855), .Z(n3812) );
  HS65_LS_NOR2X2 U14666 ( .A(n2874), .B(n2946), .Z(n3442) );
  HS65_LS_NOR2X2 U14667 ( .A(n1880), .B(n1960), .Z(n2024) );
  HS65_LS_NAND2X2 U14668 ( .A(n8787), .B(n8472), .Z(n8768) );
  HS65_LS_NAND2X2 U14669 ( .A(n8699), .B(n8412), .Z(n8680) );
  HS65_LS_NOR2X2 U14670 ( .A(n1154), .B(n1400), .Z(n1314) );
  HS65_LS_NOR2X2 U14671 ( .A(n1906), .B(n2152), .Z(n2066) );
  HS65_LS_NOR2X2 U14672 ( .A(n1129), .B(n1158), .Z(n1326) );
  HS65_LS_NOR2X2 U14673 ( .A(n1881), .B(n1910), .Z(n2078) );
  HS65_LS_NOR2X2 U14674 ( .A(n2314), .B(n2257), .Z(n2387) );
  HS65_LS_NOR2X2 U14675 ( .A(n1562), .B(n1505), .Z(n1635) );
  HS65_LS_NOR2X2 U14676 ( .A(n1186), .B(n1129), .Z(n1259) );
  HS65_LS_NOR2X2 U14677 ( .A(n1938), .B(n1881), .Z(n2011) );
  HS65_LS_NOR2X2 U14678 ( .A(n2849), .B(n3007), .Z(n3859) );
  HS65_LS_NOR2X2 U14679 ( .A(n7761), .B(n8095), .Z(n8029) );
  HS65_LS_NOR2X2 U14680 ( .A(n3003), .B(n3983), .Z(n3847) );
  HS65_LS_NOR2X2 U14681 ( .A(n1531), .B(n1549), .Z(n1662) );
  HS65_LS_NOR2X2 U14682 ( .A(n2283), .B(n2301), .Z(n2414) );
  HS65_LS_NOR2X2 U14683 ( .A(n8332), .B(n8070), .Z(n8535) );
  HS65_LS_CBI4I1X3 U14684 ( .A(n7632), .B(n7697), .C(n7639), .D(n7698), .Z(
        n7696) );
  HS65_LS_CBI4I1X3 U14685 ( .A(n7660), .B(n7735), .C(n7667), .D(n7736), .Z(
        n7734) );
  HS65_LS_NOR2X2 U14686 ( .A(n3100), .B(n2877), .Z(n3501) );
  HS65_LS_NOR2X2 U14687 ( .A(n2894), .B(n2989), .Z(n3742) );
  HS65_LS_NOR2X2 U14688 ( .A(n3043), .B(n3625), .Z(n3626) );
  HS65_LS_NOR2X2 U14689 ( .A(n7959), .B(n8361), .Z(n8071) );
  HS65_LS_NOR2X2 U14690 ( .A(n6487), .B(n6065), .Z(n6907) );
  HS65_LS_NOR2X2 U14691 ( .A(n4894), .B(n4472), .Z(n5315) );
  HS65_LS_NOR2X2 U14692 ( .A(n5008), .B(n4518), .Z(n5430) );
  HS65_LS_NOR2X2 U14693 ( .A(n6601), .B(n6111), .Z(n7022) );
  HS65_LS_NOR2X2 U14694 ( .A(n4880), .B(n4533), .Z(n5199) );
  HS65_LS_NOR2X2 U14695 ( .A(n6473), .B(n6126), .Z(n6791) );
  HS65_LS_NOR2X2 U14696 ( .A(n1155), .B(n1173), .Z(n1286) );
  HS65_LS_NOR2X2 U14697 ( .A(n8186), .B(n7661), .Z(n8836) );
  HS65_LS_NOR2X2 U14698 ( .A(n8154), .B(n7633), .Z(n8748) );
  HS65_LS_NOR2X2 U14699 ( .A(n3297), .B(n3236), .Z(n3661) );
  HS65_LS_NOR2X2 U14700 ( .A(n8164), .B(n8436), .Z(n7703) );
  HS65_LS_NOR2X2 U14701 ( .A(n8196), .B(n8447), .Z(n7741) );
  HS65_LS_NOR2X2 U14702 ( .A(n2986), .B(n3148), .Z(n3686) );
  HS65_LS_NOR2X2 U14703 ( .A(n2440), .B(n2528), .Z(n2386) );
  HS65_LS_NOR2X2 U14704 ( .A(n1688), .B(n1776), .Z(n1634) );
  HS65_LS_NOR2X2 U14705 ( .A(n2284), .B(n2328), .Z(n2479) );
  HS65_LS_NOR2X2 U14706 ( .A(n1532), .B(n1576), .Z(n1727) );
  HS65_LS_NOR2X2 U14707 ( .A(n1907), .B(n1925), .Z(n2038) );
  HS65_LS_NOR2X2 U14708 ( .A(n2371), .B(n2529), .Z(n2355) );
  HS65_LS_NOR2X2 U14709 ( .A(n1619), .B(n1777), .Z(n1603) );
  HS65_LS_NOR2X2 U14710 ( .A(n7998), .B(n8119), .Z(n8304) );
  HS65_LS_NOR2X2 U14711 ( .A(n3004), .B(n3189), .Z(n3803) );
  HS65_LS_NOR2X2 U14712 ( .A(n1312), .B(n1400), .Z(n1258) );
  HS65_LS_NOR2X2 U14713 ( .A(n2064), .B(n2152), .Z(n2010) );
  HS65_LS_NOR2X2 U14714 ( .A(n7642), .B(n7645), .Z(n8698) );
  HS65_LS_NOR2X2 U14715 ( .A(n8136), .B(n8663), .Z(n8305) );
  HS65_LS_NOR2X2 U14716 ( .A(n7670), .B(n7673), .Z(n8786) );
  HS65_LS_NOR2X2 U14717 ( .A(n1243), .B(n1401), .Z(n1227) );
  HS65_LS_NOR2X2 U14718 ( .A(n1995), .B(n2153), .Z(n1979) );
  HS65_LS_NOR2X2 U14719 ( .A(n1156), .B(n1200), .Z(n1351) );
  HS65_LS_NOR2X2 U14720 ( .A(n1908), .B(n1952), .Z(n2103) );
  HS65_LS_NOR2X2 U14721 ( .A(n3845), .B(n3983), .Z(n3406) );
  HS65_LS_NOR2X2 U14722 ( .A(n3101), .B(n2972), .Z(n3084) );
  HS65_LS_NOR2AX3 U14723 ( .A(n7709), .B(n7645), .Z(n7707) );
  HS65_LS_NOR2AX3 U14724 ( .A(n7747), .B(n7673), .Z(n7745) );
  HS65_LS_NOR2X2 U14725 ( .A(n3893), .B(n3895), .Z(n3814) );
  HS65_LS_NOR2X2 U14726 ( .A(n3263), .B(n3053), .Z(n3567) );
  HS65_LS_NOR2X2 U14727 ( .A(n3005), .B(n3208), .Z(n3884) );
  HS65_LS_NOR2X2 U14728 ( .A(n7842), .B(n7642), .Z(n8427) );
  HS65_LS_NOR2X2 U14729 ( .A(n7881), .B(n7670), .Z(n8487) );
  HS65_LS_NOR4ABX2 U14730 ( .A(n1368), .B(n1369), .C(n1370), .D(n1371), .Z(
        n1215) );
  HS65_LS_NOR3X1 U14731 ( .A(n1379), .B(n1380), .C(n1381), .Z(n1369) );
  HS65_LS_OAI212X3 U14732 ( .A(n1375), .B(n1376), .C(n1377), .D(n1186), .E(
        n1378), .Z(n1370) );
  HS65_LS_NAND4ABX3 U14733 ( .A(n1372), .B(n1138), .C(n1373), .D(n1374), .Z(
        n1371) );
  HS65_LS_NOR4ABX2 U14734 ( .A(n2496), .B(n2497), .C(n2498), .D(n2499), .Z(
        n2343) );
  HS65_LS_NOR3X1 U14735 ( .A(n2507), .B(n2508), .C(n2509), .Z(n2497) );
  HS65_LS_OAI212X3 U14736 ( .A(n2503), .B(n2504), .C(n2505), .D(n2314), .E(
        n2506), .Z(n2498) );
  HS65_LS_AOI222X2 U14737 ( .A(n901), .B(n923), .C(n899), .D(n2326), .E(n930), 
        .F(n909), .Z(n2496) );
  HS65_LS_NOR4ABX2 U14738 ( .A(n2120), .B(n2121), .C(n2122), .D(n2123), .Z(
        n1967) );
  HS65_LS_NOR3X1 U14739 ( .A(n2131), .B(n2132), .C(n2133), .Z(n2121) );
  HS65_LS_OAI212X3 U14740 ( .A(n2127), .B(n2128), .C(n2129), .D(n1938), .E(
        n2130), .Z(n2122) );
  HS65_LS_NAND4ABX3 U14741 ( .A(n2124), .B(n1890), .C(n2125), .D(n2126), .Z(
        n2123) );
  HS65_LS_NOR4ABX2 U14742 ( .A(n1744), .B(n1745), .C(n1746), .D(n1747), .Z(
        n1591) );
  HS65_LS_NOR3X1 U14743 ( .A(n1755), .B(n1756), .C(n1757), .Z(n1745) );
  HS65_LS_OAI212X3 U14744 ( .A(n1751), .B(n1752), .C(n1753), .D(n1562), .E(
        n1754), .Z(n1746) );
  HS65_LS_AOI222X2 U14745 ( .A(n819), .B(n841), .C(n817), .D(n1574), .E(n848), 
        .F(n827), .Z(n1744) );
  HS65_LS_NOR2X2 U14746 ( .A(n7817), .B(n7645), .Z(n8158) );
  HS65_LS_NOR2X2 U14747 ( .A(n7880), .B(n7673), .Z(n8190) );
  HS65_LS_NOR2X2 U14748 ( .A(n2928), .B(n3585), .Z(n3572) );
  HS65_LS_NOR2X2 U14749 ( .A(n7761), .B(n8315), .Z(n8219) );
  HS65_LS_NOR2X2 U14750 ( .A(n8136), .B(n8031), .Z(n8320) );
  HS65_LS_NAND2X2 U14751 ( .A(n7779), .B(n8379), .Z(n8333) );
  HS65_LS_NOR2X2 U14752 ( .A(n4720), .B(n4561), .Z(n5113) );
  HS65_LS_NOR2X2 U14753 ( .A(n6313), .B(n6154), .Z(n6706) );
  HS65_LS_NOR2X2 U14754 ( .A(n3625), .B(n4002), .Z(n3288) );
  HS65_LS_NAND2X2 U14755 ( .A(n7978), .B(n8436), .Z(n7852) );
  HS65_LS_NAND2X2 U14756 ( .A(n7991), .B(n8447), .Z(n7891) );
  HS65_LS_NOR2X2 U14757 ( .A(n3599), .B(n3236), .Z(n3642) );
  HS65_LS_NAND4ABX3 U14758 ( .A(n7691), .B(n7692), .C(n7693), .D(n7694), .Z(
        n7631) );
  HS65_LS_AOI212X2 U14759 ( .A(n622), .B(n7695), .C(n596), .D(n625), .E(n7696), 
        .Z(n7694) );
  HS65_LS_NAND3AX3 U14760 ( .A(n7703), .B(n7704), .C(n7705), .Z(n7692) );
  HS65_LS_MX41X4 U14761 ( .D0(n599), .S0(n620), .D1(n593), .S1(n616), .D2(n623), .S2(n584), .D3(n613), .S3(n7709), .Z(n7691) );
  HS65_LS_NAND4ABX3 U14762 ( .A(n7729), .B(n7730), .C(n7731), .D(n7732), .Z(
        n7659) );
  HS65_LS_AOI212X2 U14763 ( .A(n135), .B(n7733), .C(n109), .D(n138), .E(n7734), 
        .Z(n7732) );
  HS65_LS_NAND3AX3 U14764 ( .A(n7741), .B(n7742), .C(n7743), .Z(n7730) );
  HS65_LS_MX41X4 U14765 ( .D0(n112), .S0(n133), .D1(n106), .S1(n129), .D2(n136), .S2(n97), .D3(n126), .S3(n7747), .Z(n7729) );
  HS65_LS_NOR2X2 U14766 ( .A(n6634), .B(n7109), .Z(n6686) );
  HS65_LS_NOR2X2 U14767 ( .A(n5041), .B(n5517), .Z(n5093) );
  HS65_LS_NOR4ABX2 U14768 ( .A(n7442), .B(n7443), .C(n7444), .D(n7445), .Z(
        n7192) );
  HS65_LS_NAND3AX3 U14769 ( .A(n6906), .B(n7446), .C(n6950), .Z(n7445) );
  HS65_LS_MX41X4 U14770 ( .D0(n60), .S0(n87), .D1(n57), .S1(n89), .D2(n81), 
        .S2(n66), .D3(n84), .S3(n6184), .Z(n7444) );
  HS65_LS_AOI212X2 U14771 ( .A(n80), .B(n6921), .C(n79), .D(n58), .E(n7447), 
        .Z(n7443) );
  HS65_LS_NOR4ABX2 U14772 ( .A(n5909), .B(n5910), .C(n5911), .D(n5912), .Z(
        n5627) );
  HS65_LS_NAND3AX3 U14773 ( .A(n5429), .B(n5913), .C(n5473), .Z(n5912) );
  HS65_LS_MX41X4 U14774 ( .D0(n458), .S0(n485), .D1(n455), .S1(n487), .D2(n479), .S2(n464), .D3(n482), .S3(n4616), .Z(n5911) );
  HS65_LS_AOI212X2 U14775 ( .A(n478), .B(n5444), .C(n477), .D(n456), .E(n5914), 
        .Z(n5910) );
  HS65_LS_NOR4ABX2 U14776 ( .A(n7501), .B(n7502), .C(n7503), .D(n7504), .Z(
        n7219) );
  HS65_LS_NAND3AX3 U14777 ( .A(n7021), .B(n7505), .C(n7065), .Z(n7504) );
  HS65_LS_MX41X4 U14778 ( .D0(n281), .S0(n308), .D1(n278), .S1(n310), .D2(n302), .S2(n287), .D3(n305), .S3(n6209), .Z(n7503) );
  HS65_LS_AOI212X2 U14779 ( .A(n301), .B(n7036), .C(n300), .D(n279), .E(n7506), 
        .Z(n7502) );
  HS65_LS_NOR4ABX2 U14780 ( .A(n5850), .B(n5851), .C(n5852), .D(n5853), .Z(
        n5600) );
  HS65_LS_NAND3AX3 U14781 ( .A(n5314), .B(n5854), .C(n5358), .Z(n5853) );
  HS65_LS_MX41X4 U14782 ( .D0(n239), .S0(n266), .D1(n236), .S1(n268), .D2(n260), .S2(n245), .D3(n263), .S3(n4591), .Z(n5852) );
  HS65_LS_AOI212X2 U14783 ( .A(n259), .B(n5329), .C(n258), .D(n237), .E(n5855), 
        .Z(n5851) );
  HS65_LS_NOR4ABX2 U14784 ( .A(n5691), .B(n5692), .C(n5693), .D(n5694), .Z(
        n5583) );
  HS65_LS_NAND3AX3 U14785 ( .A(n5198), .B(n5695), .C(n5243), .Z(n5694) );
  HS65_LS_MX41X4 U14786 ( .D0(n683), .S0(n707), .D1(n689), .S1(n704), .D2(n693), .S2(n680), .D3(n702), .S3(n4531), .Z(n5693) );
  HS65_LS_AOI212X2 U14787 ( .A(n697), .B(n5213), .C(n696), .D(n690), .E(n5696), 
        .Z(n5692) );
  HS65_LS_NOR4ABX2 U14788 ( .A(n7283), .B(n7284), .C(n7285), .D(n7286), .Z(
        n7175) );
  HS65_LS_NAND3AX3 U14789 ( .A(n6790), .B(n7287), .C(n6835), .Z(n7286) );
  HS65_LS_MX41X4 U14790 ( .D0(n501), .S0(n525), .D1(n507), .S1(n522), .D2(n511), .S2(n498), .D3(n520), .S3(n6124), .Z(n7285) );
  HS65_LS_AOI212X2 U14791 ( .A(n515), .B(n6805), .C(n514), .D(n508), .E(n7288), 
        .Z(n7284) );
  HS65_LS_NOR4ABX2 U14792 ( .A(n7253), .B(n7254), .C(n7255), .D(n7256), .Z(
        n7110) );
  HS65_LS_NAND3AX3 U14793 ( .A(n6669), .B(n7257), .C(n6700), .Z(n7256) );
  HS65_LS_MX41X4 U14794 ( .D0(n544), .S0(n569), .D1(n566), .S1(n551), .D2(n541), .S2(n555), .D3(n564), .S3(n6084), .Z(n7255) );
  HS65_LS_AOI212X2 U14795 ( .A(n559), .B(n6684), .C(n558), .D(n552), .E(n7258), 
        .Z(n7254) );
  HS65_LS_NOR4ABX2 U14796 ( .A(n5661), .B(n5662), .C(n5663), .D(n5664), .Z(
        n5518) );
  HS65_LS_NAND3AX3 U14797 ( .A(n5076), .B(n5665), .C(n5107), .Z(n5664) );
  HS65_LS_MX41X4 U14798 ( .D0(n18), .S0(n43), .D1(n40), .S1(n25), .D2(n15), 
        .S2(n29), .D3(n38), .S3(n4491), .Z(n5663) );
  HS65_LS_AOI212X2 U14799 ( .A(n33), .B(n5091), .C(n32), .D(n26), .E(n5666), 
        .Z(n5662) );
  HS65_LS_CBI4I1X3 U14800 ( .A(n6153), .B(n6080), .C(n6262), .D(n6305), .Z(
        n7258) );
  HS65_LS_CBI4I1X3 U14801 ( .A(n4560), .B(n4487), .C(n4669), .D(n4712), .Z(
        n5666) );
  HS65_LS_NOR2X2 U14802 ( .A(n4989), .B(n4784), .Z(n5479) );
  HS65_LS_NOR2X2 U14803 ( .A(n4935), .B(n4745), .Z(n5364) );
  HS65_LS_NOR2X2 U14804 ( .A(n6582), .B(n6377), .Z(n7071) );
  HS65_LS_NOR2X2 U14805 ( .A(n4859), .B(n4638), .Z(n5249) );
  HS65_LS_NOR2X2 U14806 ( .A(n6452), .B(n6231), .Z(n6841) );
  HS65_LS_NOR2X2 U14807 ( .A(n6528), .B(n6338), .Z(n6956) );
  HS65_LS_NAND2X2 U14808 ( .A(n3985), .B(n3005), .Z(n2861) );
  HS65_LS_NOR2X2 U14809 ( .A(n3297), .B(n3066), .Z(n3577) );
  HS65_LS_NOR2X2 U14810 ( .A(n3263), .B(n3065), .Z(n3041) );
  HS65_LS_NOR2X2 U14811 ( .A(n8159), .B(n7833), .Z(n7683) );
  HS65_LS_NOR2X2 U14812 ( .A(n8191), .B(n7932), .Z(n7721) );
  HS65_LS_NOR2X2 U14813 ( .A(n3214), .B(n3203), .Z(n3790) );
  HS65_LS_NOR2X2 U14814 ( .A(n4495), .B(n4582), .Z(n5065) );
  HS65_LS_NOR2X2 U14815 ( .A(n6088), .B(n6175), .Z(n6658) );
  HS65_LS_NAND2X2 U14816 ( .A(n7118), .B(n7084), .Z(n6684) );
  HS65_LS_NAND2X2 U14817 ( .A(n5526), .B(n5492), .Z(n5091) );
  HS65_LS_NOR2X2 U14818 ( .A(n3470), .B(n2971), .Z(n3508) );
  HS65_LS_NAND2X2 U14819 ( .A(n7210), .B(n6064), .Z(n6921) );
  HS65_LS_NAND2X2 U14820 ( .A(n5618), .B(n4471), .Z(n5329) );
  HS65_LS_NAND2X2 U14821 ( .A(n5645), .B(n4517), .Z(n5444) );
  HS65_LS_NAND2X2 U14822 ( .A(n7237), .B(n6110), .Z(n7036) );
  HS65_LS_NAND2X2 U14823 ( .A(n5591), .B(n5508), .Z(n5213) );
  HS65_LS_NAND2X2 U14824 ( .A(n7183), .B(n7100), .Z(n6805) );
  HS65_LS_NAND2X2 U14825 ( .A(n3964), .B(n2987), .Z(n2906) );
  HS65_LS_NAND2X2 U14826 ( .A(n3942), .B(n2875), .Z(n3911) );
  HS65_LS_NAND2X2 U14827 ( .A(n3057), .B(n3282), .Z(n3247) );
  HS65_LS_NOR2X2 U14828 ( .A(n3486), .B(n2971), .Z(n3488) );
  HS65_LS_NOR2X2 U14829 ( .A(n3905), .B(n2971), .Z(n3504) );
  HS65_LS_NOR2X2 U14830 ( .A(n2943), .B(n3102), .Z(n3480) );
  HS65_LS_NAND2X2 U14831 ( .A(n1404), .B(n1156), .Z(n1141) );
  HS65_LS_NAND2X2 U14832 ( .A(n1780), .B(n1532), .Z(n1517) );
  HS65_LS_NAND2X2 U14833 ( .A(n2532), .B(n2284), .Z(n2269) );
  HS65_LS_NAND2X2 U14834 ( .A(n2156), .B(n1908), .Z(n1893) );
  HS65_LS_NOR2X2 U14835 ( .A(n5516), .B(n5026), .Z(n4689) );
  HS65_LS_NOR2X2 U14836 ( .A(n7108), .B(n6619), .Z(n6282) );
  HS65_LS_NAND2X2 U14837 ( .A(n2328), .B(n2263), .Z(n2356) );
  HS65_LS_NAND2X2 U14838 ( .A(n1576), .B(n1511), .Z(n1604) );
  HS65_LS_NOR2X2 U14839 ( .A(n6269), .B(n6086), .Z(n6670) );
  HS65_LS_NOR2X2 U14840 ( .A(n4676), .B(n4493), .Z(n5077) );
  HS65_LS_NOR2X2 U14841 ( .A(n7959), .B(n8041), .Z(n8589) );
  HS65_LS_NOR2X2 U14842 ( .A(n7862), .B(n8009), .Z(n8319) );
  HS65_LS_NOR2X2 U14843 ( .A(n8045), .B(n7954), .Z(n8565) );
  HS65_LS_NAND2X2 U14844 ( .A(n3204), .B(n3985), .Z(n3827) );
  HS65_LS_NOR2X2 U14845 ( .A(n4577), .B(n4680), .Z(n5057) );
  HS65_LS_NOR2X2 U14846 ( .A(n6170), .B(n6273), .Z(n6650) );
  HS65_LS_NOR2X2 U14847 ( .A(n3263), .B(n4103), .Z(n3269) );
  HS65_LS_NOR2X2 U14848 ( .A(n7832), .B(n7847), .Z(n7682) );
  HS65_LS_NOR2X2 U14849 ( .A(n7931), .B(n7886), .Z(n7720) );
  HS65_LS_NAND2X2 U14850 ( .A(n1200), .B(n1135), .Z(n1228) );
  HS65_LS_NAND2X2 U14851 ( .A(n1952), .B(n1887), .Z(n1980) );
  HS65_LS_NOR2X2 U14852 ( .A(n2923), .B(n3262), .Z(n3038) );
  HS65_LS_NOR2X2 U14853 ( .A(n7663), .B(n7670), .Z(n8827) );
  HS65_LS_NOR2X2 U14854 ( .A(n7635), .B(n7642), .Z(n8739) );
  HS65_LS_NOR2X2 U14855 ( .A(n3043), .B(n3282), .Z(n3647) );
  HS65_LS_NOR2X2 U14856 ( .A(n2848), .B(n3215), .Z(n3899) );
  HS65_LS_NOR2X2 U14857 ( .A(n8069), .B(n7954), .Z(n8068) );
  HS65_LS_NOR2X2 U14858 ( .A(n4509), .B(n5008), .Z(n5380) );
  HS65_LS_NOR2X2 U14859 ( .A(n4463), .B(n4894), .Z(n5265) );
  HS65_LS_NOR2X2 U14860 ( .A(n6102), .B(n6601), .Z(n6972) );
  HS65_LS_NOR2X2 U14861 ( .A(n4862), .B(n4880), .Z(n5147) );
  HS65_LS_NOR2X2 U14862 ( .A(n6455), .B(n6473), .Z(n6739) );
  HS65_LS_NOR2X2 U14863 ( .A(n6056), .B(n6487), .Z(n6857) );
  HS65_LS_NOR2X2 U14864 ( .A(n3282), .B(n3585), .Z(n3581) );
  HS65_LS_NOR2X2 U14865 ( .A(n7857), .B(n8095), .Z(n8088) );
  HS65_LS_CBI4I1X3 U14866 ( .A(n6058), .B(n6194), .C(n6481), .D(n6521), .Z(
        n7447) );
  HS65_LS_CBI4I1X3 U14867 ( .A(n4511), .B(n4613), .C(n5002), .D(n4982), .Z(
        n5914) );
  HS65_LS_CBI4I1X3 U14868 ( .A(n6104), .B(n6206), .C(n6595), .D(n6575), .Z(
        n7506) );
  HS65_LS_CBI4I1X3 U14869 ( .A(n4465), .B(n4601), .C(n4888), .D(n4928), .Z(
        n5855) );
  HS65_LS_CBI4I1X3 U14870 ( .A(n4636), .B(n4543), .C(n4874), .D(n4852), .Z(
        n5696) );
  HS65_LS_CBI4I1X3 U14871 ( .A(n6229), .B(n6136), .C(n6467), .D(n6445), .Z(
        n7288) );
  HS65_LS_NOR4ABX2 U14872 ( .A(n8145), .B(n8146), .C(n8147), .D(n8148), .Z(
        n7973) );
  HS65_LS_NOR3X1 U14873 ( .A(n7683), .B(n8157), .C(n8158), .Z(n8145) );
  HS65_LS_OAI212X3 U14874 ( .A(n7632), .B(n8149), .C(n8150), .D(n7646), .E(
        n8151), .Z(n8148) );
  HS65_LS_NAND3AX3 U14875 ( .A(n7823), .B(n8152), .C(n8153), .Z(n8147) );
  HS65_LS_NOR4ABX2 U14876 ( .A(n8177), .B(n8178), .C(n8179), .D(n8180), .Z(
        n7986) );
  HS65_LS_NOR3X1 U14877 ( .A(n7721), .B(n8189), .C(n8190), .Z(n8177) );
  HS65_LS_OAI212X3 U14878 ( .A(n7660), .B(n8181), .C(n8182), .D(n7674), .E(
        n8183), .Z(n8180) );
  HS65_LS_NAND3AX3 U14879 ( .A(n7922), .B(n8184), .C(n8185), .Z(n8179) );
  HS65_LS_NOR2X2 U14880 ( .A(n4695), .B(n4562), .Z(n5070) );
  HS65_LS_NOR2X2 U14881 ( .A(n6288), .B(n6155), .Z(n6663) );
  HS65_LS_NOR2X2 U14882 ( .A(n7871), .B(n8252), .Z(n8287) );
  HS65_LS_NOR2X2 U14883 ( .A(n3215), .B(n3208), .Z(n3824) );
  HS65_LS_NAND2X2 U14884 ( .A(n4103), .B(n2925), .Z(n3921) );
  HS65_LS_NOR2X2 U14885 ( .A(n3173), .B(n3162), .Z(n3673) );
  HS65_LS_NOR2X2 U14886 ( .A(n3058), .B(n3297), .Z(n3627) );
  HS65_LS_NOR2X2 U14887 ( .A(n7857), .B(n7999), .Z(n8286) );
  HS65_LS_NOR2X2 U14888 ( .A(n7137), .B(n6188), .Z(n6498) );
  HS65_LS_NOR2X2 U14889 ( .A(n7158), .B(n6213), .Z(n6552) );
  HS65_LS_NOR2X2 U14890 ( .A(n5545), .B(n4595), .Z(n4905) );
  HS65_LS_NOR2X2 U14891 ( .A(n5566), .B(n4620), .Z(n4959) );
  HS65_LS_NOR2X2 U14892 ( .A(n5581), .B(n5148), .Z(n4828) );
  HS65_LS_NOR2X2 U14893 ( .A(n7173), .B(n6740), .Z(n6421) );
  HS65_LS_NOR2X2 U14894 ( .A(n3728), .B(n3173), .Z(n3730) );
  HS65_LS_NAND4ABX3 U14895 ( .A(n8634), .B(n8635), .C(n8636), .D(n8637), .Z(
        n7782) );
  HS65_LS_OAI222X2 U14896 ( .A(n8326), .B(n8556), .C(n8571), .D(n7961), .E(
        n7779), .F(n8525), .Z(n8634) );
  HS65_LS_NOR3AX2 U14897 ( .A(n8515), .B(n8567), .C(n8609), .Z(n8636) );
  HS65_LS_NAND4ABX3 U14898 ( .A(n8073), .B(n8360), .C(n8622), .D(n8583), .Z(
        n8635) );
  HS65_LS_NOR2X2 U14899 ( .A(n3297), .B(n3290), .Z(n3578) );
  HS65_LS_NAND4ABX3 U14900 ( .A(n8666), .B(n8667), .C(n8668), .D(n8669), .Z(
        n7765) );
  HS65_LS_OAI222X2 U14901 ( .A(n8130), .B(n8252), .C(n8267), .D(n7859), .E(
        n7762), .F(n8220), .Z(n8666) );
  HS65_LS_NAND4ABX3 U14902 ( .A(n8028), .B(n8238), .C(n8116), .D(n8279), .Z(
        n8667) );
  HS65_LS_NOR3AX2 U14903 ( .A(n8211), .B(n8264), .C(n8305), .Z(n8668) );
  HS65_LS_NOR2X2 U14904 ( .A(n3044), .B(n2927), .Z(n3604) );
  HS65_LS_NOR2X2 U14905 ( .A(n8379), .B(n7960), .Z(n8614) );
  HS65_LS_NOR2X2 U14906 ( .A(n6064), .B(n7191), .Z(n6935) );
  HS65_LS_NOR2X2 U14907 ( .A(n4471), .B(n5599), .Z(n5343) );
  HS65_LS_NOR2X2 U14908 ( .A(n4517), .B(n5626), .Z(n5458) );
  HS65_LS_NOR2X2 U14909 ( .A(n6110), .B(n7218), .Z(n7050) );
  HS65_LS_NOR2X2 U14910 ( .A(n7100), .B(n7174), .Z(n6819) );
  HS65_LS_NOR2X2 U14911 ( .A(n5508), .B(n5582), .Z(n5227) );
  HS65_LS_NOR2X2 U14912 ( .A(n3187), .B(n2841), .Z(n3390) );
  HS65_LS_NOR2X2 U14913 ( .A(n3146), .B(n2886), .Z(n3328) );
  HS65_LS_NOR2X2 U14914 ( .A(n4559), .B(n4680), .Z(n4717) );
  HS65_LS_NOR2X2 U14915 ( .A(n6152), .B(n6273), .Z(n6310) );
  HS65_LS_NOR2X2 U14916 ( .A(n2854), .B(n3214), .Z(n3866) );
  HS65_LS_NOR2X2 U14917 ( .A(n2855), .B(n3214), .Z(n3862) );
  HS65_LS_NOR2X2 U14918 ( .A(n7964), .B(n8639), .Z(n8064) );
  HS65_LS_NOR2X2 U14919 ( .A(n1512), .B(n1530), .Z(n1620) );
  HS65_LS_NOR2X2 U14920 ( .A(n2264), .B(n2282), .Z(n2372) );
  HS65_LS_NOR4ABX2 U14921 ( .A(n6148), .B(n6149), .C(n6150), .D(n6151), .Z(
        n6077) );
  HS65_LS_NOR3X1 U14922 ( .A(n6165), .B(n6166), .C(n6167), .Z(n6148) );
  HS65_LS_OAI212X3 U14923 ( .A(n6152), .B(n6153), .C(n6154), .D(n6155), .E(
        n6156), .Z(n6151) );
  HS65_LS_NAND4ABX3 U14924 ( .A(n6157), .B(n6158), .C(n6159), .D(n6160), .Z(
        n6150) );
  HS65_LS_NOR4ABX2 U14925 ( .A(n4555), .B(n4556), .C(n4557), .D(n4558), .Z(
        n4484) );
  HS65_LS_NOR3X1 U14926 ( .A(n4572), .B(n4573), .C(n4574), .Z(n4555) );
  HS65_LS_OAI212X3 U14927 ( .A(n4559), .B(n4560), .C(n4561), .D(n4562), .E(
        n4563), .Z(n4558) );
  HS65_LS_NAND4ABX3 U14928 ( .A(n4564), .B(n4565), .C(n4566), .D(n4567), .Z(
        n4557) );
  HS65_LS_NAND2X2 U14929 ( .A(n8315), .B(n7859), .Z(n8123) );
  HS65_LS_NOR2X2 U14930 ( .A(n7778), .B(n8639), .Z(n8572) );
  HS65_LS_NOR4ABX2 U14931 ( .A(n8930), .B(n8931), .C(n8932), .D(n8933), .Z(
        n8859) );
  HS65_LS_OAI222X2 U14932 ( .A(n8639), .B(n8525), .C(n7954), .D(n7960), .E(
        n8070), .F(n8046), .Z(n8933) );
  HS65_LS_NOR3X1 U14933 ( .A(n8068), .B(n8598), .C(n8619), .Z(n8930) );
  HS65_LS_OAI212X3 U14934 ( .A(n8543), .B(n7777), .C(n7961), .D(n8069), .E(
        n8937), .Z(n8932) );
  HS65_LS_NOR2X2 U14935 ( .A(n5039), .B(n4721), .Z(n4564) );
  HS65_LS_NOR2X2 U14936 ( .A(n6632), .B(n6314), .Z(n6157) );
  HS65_LS_NOR2X2 U14937 ( .A(n5393), .B(n4990), .Z(n4787) );
  HS65_LS_NOR2X2 U14938 ( .A(n5278), .B(n4936), .Z(n4748) );
  HS65_LS_NOR2X2 U14939 ( .A(n5161), .B(n4861), .Z(n4641) );
  HS65_LS_NOR2X2 U14940 ( .A(n6985), .B(n6583), .Z(n6380) );
  HS65_LS_NOR2X2 U14941 ( .A(n6870), .B(n6529), .Z(n6341) );
  HS65_LS_NOR2X2 U14942 ( .A(n6753), .B(n6454), .Z(n6234) );
  HS65_LS_NOR2X2 U14943 ( .A(n8542), .B(n7964), .Z(n8624) );
  HS65_LS_NOR2X2 U14944 ( .A(n2299), .B(n2249), .Z(n2370) );
  HS65_LS_NOR2X2 U14945 ( .A(n1547), .B(n1497), .Z(n1618) );
  HS65_LS_NOR2X2 U14946 ( .A(n2892), .B(n3359), .Z(n3707) );
  HS65_LS_NOR2X2 U14947 ( .A(n1888), .B(n1906), .Z(n1996) );
  HS65_LS_NOR2X2 U14948 ( .A(n1136), .B(n1154), .Z(n1244) );
  HS65_LS_NOR2X2 U14949 ( .A(n1171), .B(n1214), .Z(n1307) );
  HS65_LS_NOR2X2 U14950 ( .A(n1923), .B(n1966), .Z(n2059) );
  HS65_LS_NOR2X2 U14951 ( .A(n2299), .B(n2342), .Z(n2435) );
  HS65_LS_NOR2X2 U14952 ( .A(n3102), .B(n3133), .Z(n3464) );
  HS65_LS_NOR2X2 U14953 ( .A(n1547), .B(n1590), .Z(n1683) );
  HS65_LS_NOR2X2 U14954 ( .A(n6059), .B(n6194), .Z(n6894) );
  HS65_LS_NOR2X2 U14955 ( .A(n4466), .B(n4601), .Z(n5302) );
  HS65_LS_NOR2X2 U14956 ( .A(n4512), .B(n4613), .Z(n5417) );
  HS65_LS_NOR2X2 U14957 ( .A(n6105), .B(n6206), .Z(n7009) );
  HS65_LS_NOR2X2 U14958 ( .A(n4860), .B(n4543), .Z(n5186) );
  HS65_LS_NOR2X2 U14959 ( .A(n6453), .B(n6136), .Z(n6778) );
  HS65_LS_NOR4ABX2 U14960 ( .A(n4023), .B(n4024), .C(n4025), .D(n4026), .Z(
        n3949) );
  HS65_LS_OAI222X2 U14961 ( .A(n3962), .B(n2984), .C(n3173), .D(n2986), .E(
        n3726), .F(n3147), .Z(n4026) );
  HS65_LS_NOR3X1 U14962 ( .A(n3690), .B(n3150), .C(n3330), .Z(n4023) );
  HS65_LS_OAI212X3 U14963 ( .A(n3777), .B(n2886), .C(n2987), .D(n3329), .E(
        n4027), .Z(n4025) );
  HS65_LS_NOR4ABX2 U14964 ( .A(n5519), .B(n5520), .C(n5521), .D(n5522), .Z(
        n5484) );
  HS65_LS_OAI222X2 U14965 ( .A(n5026), .B(n5523), .C(n5524), .D(n4720), .E(
        n5039), .F(n4562), .Z(n5522) );
  HS65_LS_NOR3X1 U14966 ( .A(n4570), .B(n5070), .C(n5102), .Z(n5519) );
  HS65_LS_NOR4ABX2 U14967 ( .A(n4724), .B(n4675), .C(n5042), .D(n5064), .Z(
        n5520) );
  HS65_LS_NOR4ABX2 U14968 ( .A(n7111), .B(n7112), .C(n7113), .D(n7114), .Z(
        n7076) );
  HS65_LS_OAI222X2 U14969 ( .A(n6619), .B(n7115), .C(n7116), .D(n6313), .E(
        n6632), .F(n6155), .Z(n7114) );
  HS65_LS_NOR3X1 U14970 ( .A(n6163), .B(n6663), .C(n6695), .Z(n7111) );
  HS65_LS_NOR4ABX2 U14971 ( .A(n6317), .B(n6268), .C(n6635), .D(n6657), .Z(
        n7112) );
  HS65_LS_NOR4ABX2 U14972 ( .A(n7205), .B(n7206), .C(n7207), .D(n7208), .Z(
        n7125) );
  HS65_LS_OAI222X2 U14973 ( .A(n6188), .B(n7204), .C(n7136), .D(n6528), .E(
        n6870), .F(n6339), .Z(n7208) );
  HS65_LS_NOR3X1 U14974 ( .A(n6347), .B(n6900), .C(n6945), .Z(n7205) );
  HS65_LS_OAI212X3 U14975 ( .A(n75), .B(n6051), .C(n6529), .D(n6488), .E(n7209), .Z(n7207) );
  HS65_LS_NOR4ABX2 U14976 ( .A(n7176), .B(n7177), .C(n7178), .D(n7179), .Z(
        n7092) );
  HS65_LS_OAI222X2 U14977 ( .A(n6740), .B(n7180), .C(n7181), .D(n6452), .E(
        n6753), .F(n6232), .Z(n7179) );
  HS65_LS_NOR3X1 U14978 ( .A(n6240), .B(n6784), .C(n6830), .Z(n7176) );
  HS65_LS_OAI212X3 U14979 ( .A(n516), .B(n6413), .C(n6454), .D(n6474), .E(
        n7182), .Z(n7178) );
  HS65_LS_NOR4ABX2 U14980 ( .A(n5584), .B(n5585), .C(n5586), .D(n5587), .Z(
        n5500) );
  HS65_LS_OAI222X2 U14981 ( .A(n5148), .B(n5588), .C(n5589), .D(n4859), .E(
        n5161), .F(n4639), .Z(n5587) );
  HS65_LS_NOR3X1 U14982 ( .A(n4647), .B(n5192), .C(n5238), .Z(n5584) );
  HS65_LS_OAI212X3 U14983 ( .A(n698), .B(n4820), .C(n4861), .D(n4881), .E(
        n5590), .Z(n5586) );
  HS65_LS_NOR4ABX2 U14984 ( .A(n5640), .B(n5641), .C(n5642), .D(n5643), .Z(
        n5554) );
  HS65_LS_OAI222X2 U14985 ( .A(n4620), .B(n5639), .C(n5565), .D(n4989), .E(
        n5393), .F(n4785), .Z(n5643) );
  HS65_LS_NOR3X1 U14986 ( .A(n4793), .B(n5423), .C(n5468), .Z(n5640) );
  HS65_LS_OAI212X3 U14987 ( .A(n473), .B(n4504), .C(n4990), .D(n5009), .E(
        n5644), .Z(n5642) );
  HS65_LS_NOR4ABX2 U14988 ( .A(n7232), .B(n7233), .C(n7234), .D(n7235), .Z(
        n7146) );
  HS65_LS_OAI222X2 U14989 ( .A(n6213), .B(n7231), .C(n7157), .D(n6582), .E(
        n6985), .F(n6378), .Z(n7235) );
  HS65_LS_NOR3X1 U14990 ( .A(n6386), .B(n7015), .C(n7060), .Z(n7232) );
  HS65_LS_OAI212X3 U14991 ( .A(n296), .B(n6097), .C(n6583), .D(n6602), .E(
        n7236), .Z(n7234) );
  HS65_LS_NOR4ABX2 U14992 ( .A(n5613), .B(n5614), .C(n5615), .D(n5616), .Z(
        n5533) );
  HS65_LS_OAI222X2 U14993 ( .A(n4595), .B(n5612), .C(n5544), .D(n4935), .E(
        n5278), .F(n4746), .Z(n5616) );
  HS65_LS_NOR3X1 U14994 ( .A(n4754), .B(n5308), .C(n5353), .Z(n5613) );
  HS65_LS_OAI212X3 U14995 ( .A(n254), .B(n4458), .C(n4936), .D(n4895), .E(
        n5617), .Z(n5615) );
  HS65_LS_NOR2X2 U14996 ( .A(n3187), .B(n3421), .Z(n3840) );
  HS65_LS_NOR4ABX2 U14997 ( .A(n6333), .B(n6334), .C(n6335), .D(n6336), .Z(
        n6191) );
  HS65_LS_NOR3X1 U14998 ( .A(n6349), .B(n6350), .C(n6351), .Z(n6333) );
  HS65_LS_NAND4ABX3 U14999 ( .A(n6341), .B(n6342), .C(n6343), .D(n6344), .Z(
        n6335) );
  HS65_LS_OAI212X3 U15000 ( .A(n6058), .B(n6337), .C(n6338), .D(n6339), .E(
        n6340), .Z(n6336) );
  HS65_LS_NOR4ABX2 U15001 ( .A(n4779), .B(n4780), .C(n4781), .D(n4782), .Z(
        n4610) );
  HS65_LS_NOR3X1 U15002 ( .A(n4795), .B(n4796), .C(n4797), .Z(n4779) );
  HS65_LS_NAND4ABX3 U15003 ( .A(n4787), .B(n4788), .C(n4789), .D(n4790), .Z(
        n4781) );
  HS65_LS_OAI212X3 U15004 ( .A(n4511), .B(n4783), .C(n4784), .D(n4785), .E(
        n4786), .Z(n4782) );
  HS65_LS_NOR4ABX2 U15005 ( .A(n6372), .B(n6373), .C(n6374), .D(n6375), .Z(
        n6203) );
  HS65_LS_NOR3X1 U15006 ( .A(n6388), .B(n6389), .C(n6390), .Z(n6372) );
  HS65_LS_NAND4ABX3 U15007 ( .A(n6380), .B(n6381), .C(n6382), .D(n6383), .Z(
        n6374) );
  HS65_LS_OAI212X3 U15008 ( .A(n6104), .B(n6376), .C(n6377), .D(n6378), .E(
        n6379), .Z(n6375) );
  HS65_LS_NOR4ABX2 U15009 ( .A(n4740), .B(n4741), .C(n4742), .D(n4743), .Z(
        n4598) );
  HS65_LS_NOR3X1 U15010 ( .A(n4756), .B(n4757), .C(n4758), .Z(n4740) );
  HS65_LS_NAND4ABX3 U15011 ( .A(n4748), .B(n4749), .C(n4750), .D(n4751), .Z(
        n4742) );
  HS65_LS_OAI212X3 U15012 ( .A(n4465), .B(n4744), .C(n4745), .D(n4746), .E(
        n4747), .Z(n4743) );
  HS65_LS_NOR4ABX2 U15013 ( .A(n4632), .B(n4633), .C(n4634), .D(n4635), .Z(
        n4540) );
  HS65_LS_NOR3X1 U15014 ( .A(n4649), .B(n4650), .C(n4651), .Z(n4632) );
  HS65_LS_NAND4ABX3 U15015 ( .A(n4641), .B(n4642), .C(n4643), .D(n4644), .Z(
        n4634) );
  HS65_LS_OAI212X3 U15016 ( .A(n4636), .B(n4637), .C(n4638), .D(n4639), .E(
        n4640), .Z(n4635) );
  HS65_LS_NOR4ABX2 U15017 ( .A(n6225), .B(n6226), .C(n6227), .D(n6228), .Z(
        n6133) );
  HS65_LS_NOR3X1 U15018 ( .A(n6242), .B(n6243), .C(n6244), .Z(n6225) );
  HS65_LS_NAND4ABX3 U15019 ( .A(n6234), .B(n6235), .C(n6236), .D(n6237), .Z(
        n6227) );
  HS65_LS_OAI212X3 U15020 ( .A(n6229), .B(n6230), .C(n6231), .D(n6232), .E(
        n6233), .Z(n6228) );
  HS65_LS_NOR2X2 U15021 ( .A(n8136), .B(n8018), .Z(n8264) );
  HS65_LS_NOR2X2 U15022 ( .A(n7870), .B(n8018), .Z(n8288) );
  HS65_LS_NOR2X2 U15023 ( .A(n7953), .B(n8060), .Z(n8592) );
  HS65_LS_NAND2X2 U15024 ( .A(n3893), .B(n3005), .Z(n3395) );
  HS65_LS_NOR2X2 U15025 ( .A(n1171), .B(n1121), .Z(n1242) );
  HS65_LS_NOR2X2 U15026 ( .A(n1923), .B(n1873), .Z(n1994) );
  HS65_LS_NOR2X2 U15027 ( .A(n3074), .B(n2873), .Z(n3103) );
  HS65_LS_NOR2X2 U15028 ( .A(n2944), .B(n3101), .Z(n3441) );
  HS65_LS_IVX2 U15029 ( .A(n2249), .Z(n917) );
  HS65_LS_IVX2 U15030 ( .A(n1497), .Z(n835) );
  HS65_LS_NOR2X2 U15031 ( .A(n2899), .B(n3173), .Z(n3749) );
  HS65_LS_NOR2X2 U15032 ( .A(n2900), .B(n3173), .Z(n3745) );
  HS65_LS_NOR4ABX2 U15033 ( .A(n4047), .B(n4048), .C(n4049), .D(n4050), .Z(
        n3970) );
  HS65_LS_OAI222X2 U15034 ( .A(n3983), .B(n3002), .C(n3214), .D(n3004), .E(
        n3843), .F(n3188), .Z(n4050) );
  HS65_LS_NOR3X1 U15035 ( .A(n3807), .B(n3191), .C(n3392), .Z(n4047) );
  HS65_LS_NOR4ABX2 U15036 ( .A(n3849), .B(n3420), .C(n3876), .D(n3859), .Z(
        n4048) );
  HS65_LS_NOR4ABX2 U15037 ( .A(n9039), .B(n9040), .C(n9041), .D(n9042), .Z(
        n7628) );
  HS65_LS_OAI222X2 U15038 ( .A(n7645), .B(n7832), .C(n7638), .D(n8412), .E(
        n7646), .F(n7833), .Z(n9042) );
  HS65_LS_NOR4ABX2 U15039 ( .A(n8409), .B(n8709), .C(n8433), .D(n8698), .Z(
        n9040) );
  HS65_LS_NOR3X1 U15040 ( .A(n8157), .B(n8728), .C(n8762), .Z(n9039) );
  HS65_LS_NOR4ABX2 U15041 ( .A(n9097), .B(n9098), .C(n9099), .D(n9100), .Z(
        n7656) );
  HS65_LS_OAI222X2 U15042 ( .A(n7673), .B(n7931), .C(n7666), .D(n8472), .E(
        n7674), .F(n7932), .Z(n9100) );
  HS65_LS_NOR4ABX2 U15043 ( .A(n8469), .B(n8797), .C(n8444), .D(n8786), .Z(
        n9098) );
  HS65_LS_NOR3X1 U15044 ( .A(n8189), .B(n8816), .C(n8850), .Z(n9097) );
  HS65_LS_NOR2X2 U15045 ( .A(n8003), .B(n7871), .Z(n8261) );
  HS65_LS_IVX2 U15046 ( .A(n1510), .Z(n841) );
  HS65_LS_IVX2 U15047 ( .A(n2262), .Z(n923) );
  HS65_LS_NOR2X2 U15048 ( .A(n3728), .B(n3962), .Z(n3344) );
  HS65_LS_NOR2X2 U15049 ( .A(n3845), .B(n3415), .Z(n3374) );
  HS65_LS_NOR2X2 U15050 ( .A(n3391), .B(n3415), .Z(n3398) );
  HS65_LS_NOR2X2 U15051 ( .A(n4516), .B(n4805), .Z(n5418) );
  HS65_LS_NOR2X2 U15052 ( .A(n4470), .B(n4766), .Z(n5303) );
  HS65_LS_NOR2X2 U15053 ( .A(n6109), .B(n6398), .Z(n7010) );
  HS65_LS_NOR2X2 U15054 ( .A(n4535), .B(n4659), .Z(n5187) );
  HS65_LS_NOR2X2 U15055 ( .A(n6128), .B(n6252), .Z(n6779) );
  HS65_LS_NOR2X2 U15056 ( .A(n6063), .B(n6359), .Z(n6895) );
  HS65_LS_NOR2X2 U15057 ( .A(n2850), .B(n2847), .Z(n3839) );
  HS65_LS_NOR2X2 U15058 ( .A(n7136), .B(n6529), .Z(n6347) );
  HS65_LS_NOR2X2 U15059 ( .A(n7181), .B(n6454), .Z(n6240) );
  HS65_LS_NOR2X2 U15060 ( .A(n5524), .B(n4721), .Z(n4570) );
  HS65_LS_NOR2X2 U15061 ( .A(n7116), .B(n6314), .Z(n6163) );
  HS65_LS_NOR2X2 U15062 ( .A(n5565), .B(n4990), .Z(n4793) );
  HS65_LS_NOR2X2 U15063 ( .A(n7157), .B(n6583), .Z(n6386) );
  HS65_LS_NOR2X2 U15064 ( .A(n5544), .B(n4936), .Z(n4754) );
  HS65_LS_NOR2X2 U15065 ( .A(n5589), .B(n4861), .Z(n4647) );
  HS65_LS_NOR2X2 U15066 ( .A(n2961), .B(n3133), .Z(n3498) );
  HS65_LS_NOR4ABX2 U15067 ( .A(n8982), .B(n8983), .C(n8984), .D(n8985), .Z(
        n8497) );
  HS65_LS_OAI222X2 U15068 ( .A(n8663), .B(n8220), .C(n7871), .D(n7858), .E(
        n8031), .F(n8004), .Z(n8985) );
  HS65_LS_NOR3X1 U15069 ( .A(n8026), .B(n8297), .C(n8232), .Z(n8982) );
  HS65_LS_NOR4ABX2 U15070 ( .A(n8266), .B(n8135), .C(n8124), .D(n8283), .Z(
        n8983) );
  HS65_LS_IVX2 U15071 ( .A(n1121), .Z(n876) );
  HS65_LS_IVX2 U15072 ( .A(n1873), .Z(n794) );
  HS65_LS_NOR2X2 U15073 ( .A(n2841), .B(n2849), .Z(n3198) );
  HS65_LS_NOR2X2 U15074 ( .A(n8542), .B(n7953), .Z(n8537) );
  HS65_LS_NOR2X2 U15075 ( .A(n8181), .B(n8787), .Z(n7939) );
  HS65_LS_NOR2X2 U15076 ( .A(n8149), .B(n8699), .Z(n7840) );
  HS65_LS_IVX2 U15077 ( .A(n1134), .Z(n882) );
  HS65_LS_IVX2 U15078 ( .A(n1886), .Z(n800) );
  HS65_LS_NOR2X2 U15079 ( .A(n3067), .B(n3053), .Z(n3640) );
  HS65_LS_IVX2 U15080 ( .A(n4516), .Z(n466) );
  HS65_LS_IVX2 U15081 ( .A(n4470), .Z(n247) );
  HS65_LS_IVX2 U15082 ( .A(n6109), .Z(n289) );
  HS65_LS_IVX2 U15083 ( .A(n6063), .Z(n68) );
  HS65_LS_IVX2 U15084 ( .A(n4535), .Z(n675) );
  HS65_LS_IVX2 U15085 ( .A(n6128), .Z(n493) );
  HS65_LS_NOR2X2 U15086 ( .A(n8046), .B(n7779), .Z(n8604) );
  HS65_LS_NOR2X2 U15087 ( .A(n8060), .B(n8571), .Z(n8568) );
  HS65_LS_NOR2X2 U15088 ( .A(n2856), .B(n3003), .Z(n3392) );
  HS65_LS_IVX2 U15089 ( .A(n5041), .Z(n21) );
  HS65_LS_IVX2 U15090 ( .A(n6634), .Z(n547) );
  HS65_LS_IVX2 U15091 ( .A(n4495), .Z(n10) );
  HS65_LS_IVX2 U15092 ( .A(n6088), .Z(n536) );
  HS65_LS_NOR2X2 U15093 ( .A(n3204), .B(n3421), .Z(n2857) );
  HS65_LS_NOR2X2 U15094 ( .A(n3163), .B(n3359), .Z(n2902) );
  HS65_LS_NOR4ABX2 U15095 ( .A(n3936), .B(n3937), .C(n3938), .D(n3939), .Z(
        n3907) );
  HS65_LS_OAI222X2 U15096 ( .A(n3940), .B(n3454), .C(n2971), .D(n2874), .E(
        n3484), .F(n2945), .Z(n3939) );
  HS65_LS_NOR3X1 U15097 ( .A(n3446), .B(n2948), .C(n3103), .Z(n3936) );
  HS65_LS_OAI212X3 U15098 ( .A(n3537), .B(n2973), .C(n2875), .D(n3101), .E(
        n3941), .Z(n3938) );
  HS65_LS_NAND2X2 U15099 ( .A(n3776), .B(n2987), .Z(n3333) );
  HS65_LS_NOR2X2 U15100 ( .A(n3486), .B(n3940), .Z(n3117) );
  HS65_LS_NOR2X2 U15101 ( .A(n8332), .B(n8060), .Z(n8567) );
  HS65_LS_NOR2X2 U15102 ( .A(n8060), .B(n7777), .Z(n8360) );
  HS65_LS_NOR2X2 U15103 ( .A(n4487), .B(n5516), .Z(n4583) );
  HS65_LS_NOR2X2 U15104 ( .A(n6080), .B(n7108), .Z(n6176) );
  HS65_LS_NOR2X2 U15105 ( .A(n4719), .B(n4487), .Z(n5064) );
  HS65_LS_NOR2X2 U15106 ( .A(n6312), .B(n6080), .Z(n6657) );
  HS65_LS_NOR2X2 U15107 ( .A(n7762), .B(n8136), .Z(n8246) );
  HS65_LS_NOR2X2 U15108 ( .A(n2286), .B(n2528), .Z(n2339) );
  HS65_LS_NOR2X2 U15109 ( .A(n1534), .B(n1776), .Z(n1587) );
  HS65_LS_NOR2X2 U15110 ( .A(n2283), .B(n2528), .Z(n2317) );
  HS65_LS_NOR2X2 U15111 ( .A(n1531), .B(n1776), .Z(n1565) );
  HS65_LS_NOR2X2 U15112 ( .A(n2262), .B(n2527), .Z(n2461) );
  HS65_LS_NOR2X2 U15113 ( .A(n2263), .B(n2527), .Z(n2457) );
  HS65_LS_NOR2X2 U15114 ( .A(n1511), .B(n1775), .Z(n1705) );
  HS65_LS_NOR2X2 U15115 ( .A(n1510), .B(n1775), .Z(n1709) );
  HS65_LS_IVX2 U15116 ( .A(n5395), .Z(n459) );
  HS65_LS_IVX2 U15117 ( .A(n5280), .Z(n240) );
  HS65_LS_IVX2 U15118 ( .A(n6987), .Z(n282) );
  HS65_LS_IVX2 U15119 ( .A(n5163), .Z(n685) );
  HS65_LS_IVX2 U15120 ( .A(n6755), .Z(n503) );
  HS65_LS_IVX2 U15121 ( .A(n6872), .Z(n61) );
  HS65_LS_IVX2 U15122 ( .A(n7725), .Z(n129) );
  HS65_LS_IVX2 U15123 ( .A(n7687), .Z(n616) );
  HS65_LS_NOR2X2 U15124 ( .A(n1158), .B(n1400), .Z(n1211) );
  HS65_LS_NOR2X2 U15125 ( .A(n1910), .B(n2152), .Z(n1963) );
  HS65_LS_NOR2X2 U15126 ( .A(n1155), .B(n1400), .Z(n1189) );
  HS65_LS_NOR2X2 U15127 ( .A(n1907), .B(n2152), .Z(n1941) );
  HS65_LS_NOR2X2 U15128 ( .A(n4577), .B(n4676), .Z(n5061) );
  HS65_LS_NOR2X2 U15129 ( .A(n6170), .B(n6269), .Z(n6654) );
  HS65_LS_IVX2 U15130 ( .A(n4488), .Z(n24) );
  HS65_LS_IVX2 U15131 ( .A(n6081), .Z(n550) );
  HS65_LS_NOR2X2 U15132 ( .A(n2886), .B(n2894), .Z(n3157) );
  HS65_LS_NOR2X2 U15133 ( .A(n2973), .B(n3100), .Z(n2955) );
  HS65_LS_NOR2X2 U15134 ( .A(n1135), .B(n1399), .Z(n1329) );
  HS65_LS_NOR2X2 U15135 ( .A(n1134), .B(n1399), .Z(n1333) );
  HS65_LS_NOR2X2 U15136 ( .A(n3004), .B(n3983), .Z(n3211) );
  HS65_LS_IVX2 U15137 ( .A(n4510), .Z(n454) );
  HS65_LS_IVX2 U15138 ( .A(n4464), .Z(n235) );
  HS65_LS_IVX2 U15139 ( .A(n6103), .Z(n277) );
  HS65_LS_IVX2 U15140 ( .A(n6057), .Z(n56) );
  HS65_LS_IVX2 U15141 ( .A(n4544), .Z(n688) );
  HS65_LS_IVX2 U15142 ( .A(n6137), .Z(n506) );
  HS65_LS_NOR2X2 U15143 ( .A(n3486), .B(n3127), .Z(n3083) );
  HS65_LS_NOR2X2 U15144 ( .A(n3101), .B(n3127), .Z(n3109) );
  HS65_LS_NOR2X2 U15145 ( .A(n7917), .B(n8186), .Z(n7887) );
  HS65_LS_NOR2X2 U15146 ( .A(n7818), .B(n8154), .Z(n7848) );
  HS65_LS_NOR2X2 U15147 ( .A(n2264), .B(n2342), .Z(n2475) );
  HS65_LS_NOR2X2 U15148 ( .A(n1512), .B(n1590), .Z(n1723) );
  HS65_LS_NOR2X2 U15149 ( .A(n1136), .B(n1214), .Z(n1347) );
  HS65_LS_NOR2X2 U15150 ( .A(n1888), .B(n1966), .Z(n2099) );
  HS65_LS_NOR2X2 U15151 ( .A(n7817), .B(n7847), .Z(n8433) );
  HS65_LS_NOR2X2 U15152 ( .A(n7880), .B(n7886), .Z(n8444) );
  HS65_LS_NOR2X2 U15153 ( .A(n1196), .B(n1214), .Z(n1137) );
  HS65_LS_NOR2X2 U15154 ( .A(n1948), .B(n1966), .Z(n1889) );
  HS65_LS_NOR2X2 U15155 ( .A(n2324), .B(n2342), .Z(n2265) );
  HS65_LS_NOR4ABX2 U15156 ( .A(n3974), .B(n3975), .C(n3976), .D(n3977), .Z(
        n2844) );
  HS65_LS_CBI4I1X3 U15157 ( .A(n2841), .B(n3421), .C(n3005), .D(n3384), .Z(
        n3976) );
  HS65_LS_CBI4I1X3 U15158 ( .A(n444), .B(n3215), .C(n2854), .D(n3978), .Z(
        n3977) );
  HS65_LS_NOR4ABX2 U15159 ( .A(n3797), .B(n3835), .C(n3856), .D(n3879), .Z(
        n3974) );
  HS65_LS_NOR2X2 U15160 ( .A(n1887), .B(n2151), .Z(n2081) );
  HS65_LS_NOR2X2 U15161 ( .A(n1886), .B(n2151), .Z(n2085) );
  HS65_LS_NOR2X2 U15162 ( .A(n1572), .B(n1590), .Z(n1513) );
  HS65_LS_IVX2 U15163 ( .A(n2899), .Z(n648) );
  HS65_LS_NOR3AX2 U15164 ( .A(n4067), .B(n4068), .C(n3908), .Z(n4064) );
  HS65_LS_OAI21X2 U15165 ( .A(n2965), .B(n2946), .C(n4074), .Z(n4068) );
  HS65_LS_NOR2X2 U15166 ( .A(n8018), .B(n8267), .Z(n8263) );
  HS65_LS_NOR2X2 U15167 ( .A(n7108), .B(n6269), .Z(n6711) );
  HS65_LS_NOR2X2 U15168 ( .A(n5516), .B(n4676), .Z(n5118) );
  HS65_LS_NOR2X2 U15169 ( .A(n8150), .B(n8699), .Z(n8156) );
  HS65_LS_NOR2X2 U15170 ( .A(n8182), .B(n8787), .Z(n8188) );
  HS65_LS_NOR2X2 U15171 ( .A(n6194), .B(n7204), .Z(n6484) );
  HS65_LS_NOR2X2 U15172 ( .A(n6206), .B(n7231), .Z(n6598) );
  HS65_LS_NOR2X2 U15173 ( .A(n6528), .B(n7204), .Z(n6361) );
  HS65_LS_NOR2X2 U15174 ( .A(n4989), .B(n5639), .Z(n4807) );
  HS65_LS_NOR2X2 U15175 ( .A(n6582), .B(n7231), .Z(n6400) );
  HS65_LS_NOR2X2 U15176 ( .A(n4601), .B(n5612), .Z(n4891) );
  HS65_LS_NOR2X2 U15177 ( .A(n4613), .B(n5639), .Z(n5005) );
  HS65_LS_NOR2X2 U15178 ( .A(n4935), .B(n5612), .Z(n4768) );
  HS65_LS_NOR2X2 U15179 ( .A(n4859), .B(n5588), .Z(n4661) );
  HS65_LS_NOR2X2 U15180 ( .A(n4543), .B(n5588), .Z(n4877) );
  HS65_LS_NOR2X2 U15181 ( .A(n6452), .B(n7180), .Z(n6254) );
  HS65_LS_NOR2X2 U15182 ( .A(n6136), .B(n7180), .Z(n6470) );
  HS65_LS_NOR2X2 U15183 ( .A(n8154), .B(n7687), .Z(n8730) );
  HS65_LS_NOR2X2 U15184 ( .A(n8186), .B(n7725), .Z(n8818) );
  HS65_LS_NOR2X2 U15185 ( .A(n2249), .B(n2257), .Z(n2310) );
  HS65_LS_NOR2X2 U15186 ( .A(n1121), .B(n1129), .Z(n1182) );
  HS65_LS_NOR2X2 U15187 ( .A(n1873), .B(n1881), .Z(n1934) );
  HS65_LS_NOR2X2 U15188 ( .A(n1497), .B(n1505), .Z(n1558) );
  HS65_LS_NOR2X2 U15189 ( .A(n8315), .B(n7862), .Z(n8237) );
  HS65_LS_NOR2X2 U15190 ( .A(n4504), .B(n4783), .Z(n4987) );
  HS65_LS_NOR2X2 U15191 ( .A(n4458), .B(n4744), .Z(n4933) );
  HS65_LS_NOR2X2 U15192 ( .A(n4820), .B(n4637), .Z(n4857) );
  HS65_LS_NOR2X2 U15193 ( .A(n6097), .B(n6376), .Z(n6580) );
  HS65_LS_NOR2X2 U15194 ( .A(n6413), .B(n6230), .Z(n6450) );
  HS65_LS_NOR2X2 U15195 ( .A(n6051), .B(n6337), .Z(n6526) );
  HS65_LS_NOR2X2 U15196 ( .A(n2529), .B(n2328), .Z(n2481) );
  HS65_LS_NOR2X2 U15197 ( .A(n1777), .B(n1576), .Z(n1729) );
  HS65_LS_NOR2X2 U15198 ( .A(n3043), .B(n3067), .Z(n3260) );
  HS65_LS_NOR2AX3 U15199 ( .A(n4491), .B(n4722), .Z(n5062) );
  HS65_LS_NOR2AX3 U15200 ( .A(n6084), .B(n6315), .Z(n6655) );
  HS65_LS_NOR2X2 U15201 ( .A(n7686), .B(n7818), .Z(n8715) );
  HS65_LS_NOR2X2 U15202 ( .A(n7724), .B(n7917), .Z(n8803) );
  HS65_LS_NOR2X2 U15203 ( .A(n2900), .B(n3146), .Z(n3748) );
  HS65_LS_OAI21X2 U15204 ( .A(n2973), .B(n3074), .C(n3075), .Z(n3073) );
  HS65_LS_OAI21X2 U15205 ( .A(n2841), .B(n2856), .C(n3366), .Z(n3365) );
  HS65_LS_NOR2X2 U15206 ( .A(n7832), .B(n7633), .Z(n7803) );
  HS65_LS_NOR2X2 U15207 ( .A(n7931), .B(n7661), .Z(n7903) );
  HS65_LS_NOR4ABX2 U15208 ( .A(n4196), .B(n4197), .C(n4198), .D(n4199), .Z(
        n3910) );
  HS65_LS_CBI4I1X3 U15209 ( .A(n2973), .B(n3133), .C(n2875), .D(n3093), .Z(
        n4198) );
  HS65_LS_CBI4I1X3 U15210 ( .A(n220), .B(n2972), .C(n3470), .D(n4200), .Z(
        n4199) );
  HS65_LS_NOR4ABX2 U15211 ( .A(n3436), .B(n3476), .C(n3497), .D(n3521), .Z(
        n4196) );
  HS65_LS_NOR2X2 U15212 ( .A(n2848), .B(n3893), .Z(n3802) );
  HS65_LS_NOR2X2 U15213 ( .A(n1401), .B(n1200), .Z(n1353) );
  HS65_LS_NOR2X2 U15214 ( .A(n2153), .B(n1952), .Z(n2105) );
  HS65_LS_NOR2X2 U15215 ( .A(n2263), .B(n2299), .Z(n2460) );
  HS65_LS_NOR2X2 U15216 ( .A(n1511), .B(n1547), .Z(n1708) );
  HS65_LS_NAND2X2 U15217 ( .A(n7870), .B(n8220), .Z(n7875) );
  HS65_LS_NOR2X2 U15218 ( .A(n3057), .B(n3066), .Z(n3605) );
  HS65_LS_NAND2X2 U15219 ( .A(n7955), .B(n7960), .Z(n8043) );
  HS65_LS_NOR2X2 U15220 ( .A(n8315), .B(n7870), .Z(n8310) );
  HS65_LS_NOR2X2 U15221 ( .A(n4722), .B(n4676), .Z(n5025) );
  HS65_LS_NOR2X2 U15222 ( .A(n6315), .B(n6269), .Z(n6618) );
  HS65_LS_NOR2X2 U15223 ( .A(n8160), .B(n7638), .Z(n8683) );
  HS65_LS_NOR2X2 U15224 ( .A(n8192), .B(n7666), .Z(n8771) );
  HS65_LS_NAND2X2 U15225 ( .A(n5492), .B(n5026), .Z(n4497) );
  HS65_LS_NAND2X2 U15226 ( .A(n7084), .B(n6619), .Z(n6090) );
  HS65_LS_NOR2X2 U15227 ( .A(n1135), .B(n1171), .Z(n1332) );
  HS65_LS_NOR2X2 U15228 ( .A(n8130), .B(n8267), .Z(n8103) );
  HS65_LS_NAND2X2 U15229 ( .A(n4517), .B(n4620), .Z(n4514) );
  HS65_LS_NAND2X2 U15230 ( .A(n4471), .B(n4595), .Z(n4468) );
  HS65_LS_NAND2X2 U15231 ( .A(n6110), .B(n6213), .Z(n6107) );
  HS65_LS_NAND2X2 U15232 ( .A(n5508), .B(n5148), .Z(n4537) );
  HS65_LS_NAND2X2 U15233 ( .A(n7100), .B(n6740), .Z(n6130) );
  HS65_LS_NAND2X2 U15234 ( .A(n6064), .B(n6188), .Z(n6061) );
  HS65_LS_IVX2 U15235 ( .A(n2986), .Z(n641) );
  HS65_LS_NOR2X2 U15236 ( .A(n8326), .B(n8571), .Z(n8344) );
  HS65_LS_NOR2X2 U15237 ( .A(n4680), .B(n4494), .Z(n4714) );
  HS65_LS_NOR2X2 U15238 ( .A(n6273), .B(n6087), .Z(n6307) );
  HS65_LS_NAND2X2 U15239 ( .A(n2850), .B(n3004), .Z(n3206) );
  HS65_LS_NOR2X2 U15240 ( .A(n1887), .B(n1923), .Z(n2084) );
  HS65_LS_NOR2X2 U15241 ( .A(n8030), .B(n7871), .Z(n8026) );
  HS65_LS_NOR2X2 U15242 ( .A(n2899), .B(n3726), .Z(n3699) );
  HS65_LS_NOR4ABX2 U15243 ( .A(n3953), .B(n3954), .C(n3955), .D(n3956), .Z(
        n2889) );
  HS65_LS_CBI4I1X3 U15244 ( .A(n2886), .B(n3359), .C(n2987), .D(n3322), .Z(
        n3955) );
  HS65_LS_CBI4I1X3 U15245 ( .A(n668), .B(n3174), .C(n2899), .D(n3957), .Z(
        n3956) );
  HS65_LS_NOR4ABX2 U15246 ( .A(n3680), .B(n3719), .C(n3739), .D(n3762), .Z(
        n3953) );
  HS65_LS_NOR2X2 U15247 ( .A(n8069), .B(n8051), .Z(n8345) );
  HS65_LS_NOR2X2 U15248 ( .A(n2256), .B(n2529), .Z(n2509) );
  HS65_LS_NOR2X2 U15249 ( .A(n1504), .B(n1777), .Z(n1757) );
  HS65_LS_NOR2X2 U15250 ( .A(n7632), .B(n7687), .Z(n7799) );
  HS65_LS_NOR2X2 U15251 ( .A(n7660), .B(n7725), .Z(n7899) );
  HS65_LS_NAND2X2 U15252 ( .A(n7872), .B(n7858), .Z(n8001) );
  HS65_LS_NOR2X2 U15253 ( .A(n6057), .B(n7191), .Z(n6951) );
  HS65_LS_NOR2X2 U15254 ( .A(n6103), .B(n7218), .Z(n7066) );
  HS65_LS_NOR2X2 U15255 ( .A(n4510), .B(n5626), .Z(n5474) );
  HS65_LS_NOR2X2 U15256 ( .A(n4464), .B(n5599), .Z(n5359) );
  HS65_LS_NOR2X2 U15257 ( .A(n4544), .B(n5582), .Z(n5244) );
  HS65_LS_NOR2X2 U15258 ( .A(n6137), .B(n7174), .Z(n6836) );
  HS65_LS_NOR2X2 U15259 ( .A(n2527), .B(n2328), .Z(n2433) );
  HS65_LS_NOR2X2 U15260 ( .A(n1775), .B(n1576), .Z(n1681) );
  HS65_LS_IVX2 U15261 ( .A(n8252), .Z(n369) );
  HS65_LS_IVX2 U15262 ( .A(n8556), .Z(n322) );
  HS65_LS_NOR2X2 U15263 ( .A(n3280), .B(n3297), .Z(n3579) );
  HS65_LS_NOR2X2 U15264 ( .A(n2893), .B(n3776), .Z(n3685) );
  HS65_LS_NOR2X2 U15265 ( .A(n2878), .B(n2971), .Z(n3430) );
  HS65_LS_NOR2X2 U15266 ( .A(n2901), .B(n2985), .Z(n3330) );
  HS65_LS_IVX2 U15267 ( .A(n2973), .Z(n191) );
  HS65_LS_NOR2X2 U15268 ( .A(n1128), .B(n1401), .Z(n1381) );
  HS65_LS_NOR2X2 U15269 ( .A(n1880), .B(n2153), .Z(n2133) );
  HS65_LS_CBI4I1X3 U15270 ( .A(n2336), .B(n2301), .C(n2262), .D(n2425), .Z(
        n2424) );
  HS65_LS_CBI4I1X3 U15271 ( .A(n1584), .B(n1549), .C(n1510), .D(n1673), .Z(
        n1672) );
  HS65_LS_NOR2X2 U15272 ( .A(n7686), .B(n7645), .Z(n8760) );
  HS65_LS_NOR2X2 U15273 ( .A(n7724), .B(n7673), .Z(n8848) );
  HS65_LS_NOR2X2 U15274 ( .A(n3187), .B(n3845), .Z(n3841) );
  HS65_LS_NOR2X2 U15275 ( .A(n2855), .B(n3893), .Z(n3889) );
  HS65_LS_NOR2X2 U15276 ( .A(n7959), .B(n7954), .Z(n8593) );
  HS65_LS_NOR2X2 U15277 ( .A(n1399), .B(n1200), .Z(n1305) );
  HS65_LS_NOR2X2 U15278 ( .A(n2151), .B(n1952), .Z(n2057) );
  HS65_LS_CBI4I1X3 U15279 ( .A(n1208), .B(n1173), .C(n1134), .D(n1297), .Z(
        n1296) );
  HS65_LS_NOR2X2 U15280 ( .A(n8159), .B(n7638), .Z(n8157) );
  HS65_LS_NOR2X2 U15281 ( .A(n8191), .B(n7666), .Z(n8189) );
  HS65_LS_NOR2X2 U15282 ( .A(n3263), .B(n3066), .Z(n3246) );
  HS65_LS_NOR2X2 U15283 ( .A(n1171), .B(n1312), .Z(n1308) );
  HS65_LS_NOR2X2 U15284 ( .A(n1923), .B(n2064), .Z(n2060) );
  HS65_LS_NOR2X2 U15285 ( .A(n1547), .B(n1688), .Z(n1684) );
  HS65_LS_NOR2X2 U15286 ( .A(n2299), .B(n2440), .Z(n2436) );
  HS65_LS_IVX2 U15287 ( .A(n8525), .Z(n323) );
  HS65_LS_OAI21X2 U15288 ( .A(n7760), .B(n8095), .C(n8650), .Z(n8649) );
  HS65_LS_NOR2X2 U15289 ( .A(n3625), .B(n3262), .Z(n3265) );
  HS65_LS_CBI4I1X3 U15290 ( .A(n1960), .B(n1925), .C(n1886), .D(n2049), .Z(
        n2048) );
  HS65_LS_IVX2 U15291 ( .A(n2987), .Z(n661) );
  HS65_LS_IVX2 U15292 ( .A(n3005), .Z(n437) );
  HS65_LS_IVX2 U15293 ( .A(n2875), .Z(n212) );
  HS65_LS_NOR2X2 U15294 ( .A(n4800), .B(n5008), .Z(n4519) );
  HS65_LS_NOR2X2 U15295 ( .A(n4761), .B(n4894), .Z(n4473) );
  HS65_LS_NOR2X2 U15296 ( .A(n6393), .B(n6601), .Z(n6112) );
  HS65_LS_NOR2X2 U15297 ( .A(n4654), .B(n4880), .Z(n5183) );
  HS65_LS_NOR2X2 U15298 ( .A(n6247), .B(n6473), .Z(n6775) );
  HS65_LS_NOR2X2 U15299 ( .A(n6354), .B(n6487), .Z(n6066) );
  HS65_LS_IVX2 U15300 ( .A(n3845), .Z(n411) );
  HS65_LS_NOR2AX3 U15301 ( .A(n4491), .B(n4695), .Z(n4687) );
  HS65_LS_NOR2AX3 U15302 ( .A(n6084), .B(n6288), .Z(n6280) );
  HS65_LS_CBI4I1X3 U15303 ( .A(n3353), .B(n3148), .C(n2899), .D(n3713), .Z(
        n3712) );
  HS65_LS_NOR2X2 U15304 ( .A(n3214), .B(n3208), .Z(n3838) );
  HS65_LS_IVX2 U15305 ( .A(n2314), .Z(n920) );
  HS65_LS_IVX2 U15306 ( .A(n1562), .Z(n838) );
  HS65_LS_IVX2 U15307 ( .A(n7859), .Z(n404) );
  HS65_LS_NOR2X2 U15308 ( .A(n3146), .B(n3728), .Z(n3724) );
  HS65_LS_IVX2 U15309 ( .A(n8787), .Z(n114) );
  HS65_LS_IVX2 U15310 ( .A(n8699), .Z(n601) );
  HS65_LS_NAND2X2 U15311 ( .A(n2946), .B(n2944), .Z(n2951) );
  HS65_LS_NOR2X2 U15312 ( .A(n3905), .B(n2944), .Z(n3507) );
  HS65_LS_NOR2X2 U15313 ( .A(n2855), .B(n3187), .Z(n3865) );
  HS65_LS_NAND2X2 U15314 ( .A(n7885), .B(n7931), .Z(n7883) );
  HS65_LS_NAND2X2 U15315 ( .A(n7846), .B(n7832), .Z(n7844) );
  HS65_LS_IVX2 U15316 ( .A(n2925), .Z(n166) );
  HS65_LS_NAND4ABX3 U15317 ( .A(n3339), .B(n3340), .C(n3341), .D(n3342), .Z(
        n2981) );
  HS65_LS_NOR3X1 U15318 ( .A(n3343), .B(n3344), .C(n3345), .Z(n3342) );
  HS65_LS_OAI212X3 U15319 ( .A(n3349), .B(n2887), .C(n3162), .D(n2901), .E(
        n3350), .Z(n3339) );
  HS65_LS_AOI222X2 U15320 ( .A(n643), .B(n665), .C(n646), .D(n667), .E(n644), 
        .F(n658), .Z(n3341) );
  HS65_LS_CBI4I1X3 U15321 ( .A(n7639), .B(n8150), .C(n7634), .D(n8690), .Z(
        n8689) );
  HS65_LS_CBI4I1X3 U15322 ( .A(n7667), .B(n8182), .C(n7662), .D(n8778), .Z(
        n8777) );
  HS65_LS_IVX2 U15323 ( .A(n1186), .Z(n879) );
  HS65_LS_IVX2 U15324 ( .A(n1938), .Z(n797) );
  HS65_LS_NOR2X2 U15325 ( .A(n3985), .B(n2841), .Z(n3386) );
  HS65_LS_NOR2X2 U15326 ( .A(n3964), .B(n2886), .Z(n3324) );
  HS65_LS_NOR2X2 U15327 ( .A(n6194), .B(n7137), .Z(n6360) );
  HS65_LS_NOR2X2 U15328 ( .A(n4613), .B(n5566), .Z(n4806) );
  HS65_LS_NOR2X2 U15329 ( .A(n6206), .B(n7158), .Z(n6399) );
  HS65_LS_NOR2X2 U15330 ( .A(n4601), .B(n5545), .Z(n4767) );
  HS65_LS_NOR2X2 U15331 ( .A(n4543), .B(n5581), .Z(n4660) );
  HS65_LS_NOR2X2 U15332 ( .A(n6136), .B(n7173), .Z(n6253) );
  HS65_LS_NOR2X2 U15333 ( .A(n2900), .B(n3776), .Z(n3772) );
  HS65_LS_IVX2 U15334 ( .A(n1312), .Z(n888) );
  HS65_LS_IVX2 U15335 ( .A(n2064), .Z(n806) );
  HS65_LS_IVX2 U15336 ( .A(n2440), .Z(n929) );
  HS65_LS_IVX2 U15337 ( .A(n1688), .Z(n847) );
  HS65_LS_NAND2X2 U15338 ( .A(n2301), .B(n2299), .Z(n2306) );
  HS65_LS_NAND2X2 U15339 ( .A(n1549), .B(n1547), .Z(n1554) );
  HS65_LS_NOR3X1 U15340 ( .A(n4306), .B(n2845), .C(n3973), .Z(n4303) );
  HS65_LS_OAI21X2 U15341 ( .A(n3208), .B(n3189), .C(n3979), .Z(n4306) );
  HS65_LS_NOR3X1 U15342 ( .A(n4247), .B(n2890), .C(n3952), .Z(n4244) );
  HS65_LS_OAI21X2 U15343 ( .A(n3167), .B(n3148), .C(n3958), .Z(n4247) );
  HS65_LS_NOR2X2 U15344 ( .A(n3895), .B(n2842), .Z(n3200) );
  HS65_LS_IVX2 U15345 ( .A(n7842), .Z(n612) );
  HS65_LS_IVX2 U15346 ( .A(n7881), .Z(n125) );
  HS65_LS_NOR2X2 U15347 ( .A(n7137), .B(n6487), .Z(n6932) );
  HS65_LS_NOR2X2 U15348 ( .A(n5545), .B(n4894), .Z(n5340) );
  HS65_LS_NOR2X2 U15349 ( .A(n5566), .B(n5008), .Z(n5455) );
  HS65_LS_NOR2X2 U15350 ( .A(n7158), .B(n6601), .Z(n7047) );
  HS65_LS_NOR2X2 U15351 ( .A(n7173), .B(n6473), .Z(n6816) );
  HS65_LS_NOR2X2 U15352 ( .A(n5581), .B(n4880), .Z(n5224) );
  HS65_LS_NOR2X2 U15353 ( .A(n3329), .B(n3174), .Z(n3313) );
  HS65_LS_NOR2X2 U15354 ( .A(n2532), .B(n2249), .Z(n2366) );
  HS65_LS_NOR2X2 U15355 ( .A(n1780), .B(n1497), .Z(n1614) );
  HS65_LS_NAND2X2 U15356 ( .A(n3282), .B(n3599), .Z(n2922) );
  HS65_LS_IVX2 U15357 ( .A(n3127), .Z(n226) );
  HS65_LS_NOR2X2 U15358 ( .A(n4559), .B(n5526), .Z(n4729) );
  HS65_LS_NOR2X2 U15359 ( .A(n6152), .B(n7118), .Z(n6322) );
  HS65_LS_NAND2X2 U15360 ( .A(n1173), .B(n1171), .Z(n1178) );
  HS65_LS_AOI12X2 U15361 ( .A(n2886), .B(n3728), .C(n3726), .Z(n3963) );
  HS65_LS_NOR2X2 U15362 ( .A(n6186), .B(n6051), .Z(n6523) );
  HS65_LS_NOR2X2 U15363 ( .A(n6211), .B(n6097), .Z(n6577) );
  HS65_LS_NOR2X2 U15364 ( .A(n4618), .B(n4504), .Z(n4984) );
  HS65_LS_NOR2X2 U15365 ( .A(n4593), .B(n4458), .Z(n4930) );
  HS65_LS_NOR2X2 U15366 ( .A(n4534), .B(n4820), .Z(n4854) );
  HS65_LS_NOR2X2 U15367 ( .A(n6127), .B(n6413), .Z(n6447) );
  HS65_LS_NOR2X2 U15368 ( .A(n1404), .B(n1121), .Z(n1238) );
  HS65_LS_NOR2X2 U15369 ( .A(n2156), .B(n1873), .Z(n1990) );
  HS65_LS_CBI4I1X3 U15370 ( .A(n2943), .B(n2877), .C(n3127), .D(n3444), .Z(
        n4066) );
  HS65_LS_NOR2X2 U15371 ( .A(n2878), .B(n2972), .Z(n3541) );
  HS65_LS_IVX2 U15372 ( .A(n3778), .Z(n643) );
  HS65_LS_NAND2X2 U15373 ( .A(n3148), .B(n3146), .Z(n3153) );
  HS65_LS_NOR2X2 U15374 ( .A(n1136), .B(n1158), .Z(n1248) );
  HS65_LS_NOR2X2 U15375 ( .A(n1888), .B(n1910), .Z(n2000) );
  HS65_LS_NOR2X2 U15376 ( .A(n1512), .B(n1534), .Z(n1624) );
  HS65_LS_NOR2X2 U15377 ( .A(n2264), .B(n2286), .Z(n2376) );
  HS65_LS_NOR2X2 U15378 ( .A(n4720), .B(n5523), .Z(n4584) );
  HS65_LS_NOR2X2 U15379 ( .A(n6313), .B(n7115), .Z(n6177) );
  HS65_LS_IVX2 U15380 ( .A(n3728), .Z(n634) );
  HS65_LS_IVX2 U15381 ( .A(n1511), .Z(n836) );
  HS65_LS_IVX2 U15382 ( .A(n2263), .Z(n918) );
  HS65_LS_OAI21X2 U15383 ( .A(n2886), .B(n2901), .C(n3304), .Z(n3303) );
  HS65_LS_NOR2X2 U15384 ( .A(n4487), .B(n5523), .Z(n4673) );
  HS65_LS_NOR2X2 U15385 ( .A(n6080), .B(n7115), .Z(n6266) );
  HS65_LS_NAND2X2 U15386 ( .A(n1925), .B(n1923), .Z(n1930) );
  HS65_LS_OAI21X2 U15387 ( .A(n8361), .B(n8332), .C(n8616), .Z(n8900) );
  HS65_LS_NOR2X2 U15388 ( .A(n3074), .B(n2877), .Z(n3107) );
  HS65_LS_NOR2X2 U15389 ( .A(n2856), .B(n3007), .Z(n3396) );
  HS65_LS_NOR2X2 U15390 ( .A(n2944), .B(n3470), .Z(n3455) );
  HS65_LS_NAND2X2 U15391 ( .A(n3189), .B(n3187), .Z(n3194) );
  HS65_LS_NOR2X2 U15392 ( .A(n7667), .B(n8186), .Z(n7888) );
  HS65_LS_NOR2X2 U15393 ( .A(n7639), .B(n8154), .Z(n7849) );
  HS65_LS_OAI21X2 U15394 ( .A(n2504), .B(n2335), .C(n2565), .Z(n2564) );
  HS65_LS_OAI21X2 U15395 ( .A(n917), .B(n920), .C(n901), .Z(n2565) );
  HS65_LS_OAI21X2 U15396 ( .A(n2128), .B(n1959), .C(n2189), .Z(n2188) );
  HS65_LS_OAI21X2 U15397 ( .A(n794), .B(n797), .C(n778), .Z(n2189) );
  HS65_LS_OAI21X2 U15398 ( .A(n1752), .B(n1583), .C(n1813), .Z(n1812) );
  HS65_LS_OAI21X2 U15399 ( .A(n835), .B(n838), .C(n819), .Z(n1813) );
  HS65_LS_OAI21X2 U15400 ( .A(n1376), .B(n1207), .C(n1437), .Z(n1436) );
  HS65_LS_OAI21X2 U15401 ( .A(n876), .B(n879), .C(n860), .Z(n1437) );
  HS65_LS_NOR2X2 U15402 ( .A(n3942), .B(n2973), .Z(n3095) );
  HS65_LS_NAND2X2 U15403 ( .A(n569), .B(n6084), .Z(n6690) );
  HS65_LS_NAND2X2 U15404 ( .A(n43), .B(n4491), .Z(n5097) );
  HS65_LS_NOR2X2 U15405 ( .A(n8335), .B(n8525), .Z(n7773) );
  HS65_LS_IVX2 U15406 ( .A(n1135), .Z(n877) );
  HS65_LS_IVX2 U15407 ( .A(n1887), .Z(n795) );
  HS65_LS_NOR2X2 U15408 ( .A(n7964), .B(n7954), .Z(n8517) );
  HS65_LS_AOI12X2 U15409 ( .A(n4504), .B(n5395), .C(n5393), .Z(n5569) );
  HS65_LS_AOI12X2 U15410 ( .A(n6097), .B(n6987), .C(n6985), .Z(n7161) );
  HS65_LS_AOI12X2 U15411 ( .A(n6051), .B(n6872), .C(n6870), .Z(n7140) );
  HS65_LS_AOI12X2 U15412 ( .A(n4458), .B(n5280), .C(n5278), .Z(n5548) );
  HS65_LS_NOR2X2 U15413 ( .A(n3536), .B(n3538), .Z(n3453) );
  HS65_LS_IVX2 U15414 ( .A(n2841), .Z(n425) );
  HS65_LS_IVX2 U15415 ( .A(n2886), .Z(n649) );
  HS65_LS_NOR2X2 U15416 ( .A(n2944), .B(n3486), .Z(n3481) );
  HS65_LS_NOR2X2 U15417 ( .A(n2928), .B(n3065), .Z(n3556) );
  HS65_LS_NOR2X2 U15418 ( .A(n8881), .B(n7777), .Z(n8356) );
  HS65_LS_NOR2X2 U15419 ( .A(n8671), .B(n7760), .Z(n8114) );
  HS65_LS_IVX2 U15420 ( .A(n8571), .Z(n327) );
  HS65_LS_NOR2X2 U15421 ( .A(n1376), .B(n1186), .Z(n1367) );
  HS65_LS_NOR2X2 U15422 ( .A(n2504), .B(n2314), .Z(n2495) );
  HS65_LS_NOR2X2 U15423 ( .A(n2128), .B(n1938), .Z(n2119) );
  HS65_LS_NOR2X2 U15424 ( .A(n1752), .B(n1562), .Z(n1743) );
  HS65_LS_CBI4I6X2 U15425 ( .A(n903), .B(n908), .C(n917), .D(n2321), .Z(n2319)
         );
  HS65_LS_AOI12X2 U15426 ( .A(n2262), .B(n2258), .C(n2250), .Z(n2321) );
  HS65_LS_CBI4I6X2 U15427 ( .A(n821), .B(n826), .C(n835), .D(n1569), .Z(n1567)
         );
  HS65_LS_AOI12X2 U15428 ( .A(n1510), .B(n1506), .C(n1498), .Z(n1569) );
  HS65_LS_CBI4I6X2 U15429 ( .A(n862), .B(n867), .C(n876), .D(n1193), .Z(n1191)
         );
  HS65_LS_AOI12X2 U15430 ( .A(n1134), .B(n1130), .C(n1122), .Z(n1193) );
  HS65_LS_CBI4I6X2 U15431 ( .A(n780), .B(n785), .C(n794), .D(n1945), .Z(n1943)
         );
  HS65_LS_AOI12X2 U15432 ( .A(n1886), .B(n1882), .C(n1874), .Z(n1945) );
  HS65_LS_IVX2 U15433 ( .A(n4504), .Z(n467) );
  HS65_LS_IVX2 U15434 ( .A(n4458), .Z(n248) );
  HS65_LS_IVX2 U15435 ( .A(n4820), .Z(n677) );
  HS65_LS_IVX2 U15436 ( .A(n6097), .Z(n290) );
  HS65_LS_IVX2 U15437 ( .A(n6051), .Z(n69) );
  HS65_LS_IVX2 U15438 ( .A(n6413), .Z(n495) );
  HS65_LS_NOR2X2 U15439 ( .A(n3281), .B(n3066), .Z(n3564) );
  HS65_LS_NAND2X2 U15440 ( .A(n8019), .B(n8018), .Z(n7753) );
  HS65_LS_NAND2X2 U15441 ( .A(n8061), .B(n8060), .Z(n7784) );
  HS65_LS_NAND2X2 U15442 ( .A(n2263), .B(n2281), .Z(n2260) );
  HS65_LS_NAND2X2 U15443 ( .A(n1511), .B(n1529), .Z(n1508) );
  HS65_LS_NAND2X2 U15444 ( .A(n7666), .B(n7672), .Z(n8838) );
  HS65_LS_NAND2X2 U15445 ( .A(n7638), .B(n7644), .Z(n8750) );
  HS65_LS_NAND2X2 U15446 ( .A(n87), .B(n6184), .Z(n6927) );
  HS65_LS_NAND2X2 U15447 ( .A(n266), .B(n4591), .Z(n5335) );
  HS65_LS_NAND2X2 U15448 ( .A(n485), .B(n4616), .Z(n5450) );
  HS65_LS_NAND2X2 U15449 ( .A(n308), .B(n6209), .Z(n7042) );
  HS65_LS_NAND2X2 U15450 ( .A(n525), .B(n6124), .Z(n6811) );
  HS65_LS_NAND2X2 U15451 ( .A(n707), .B(n4531), .Z(n5219) );
  HS65_LS_NAND2X2 U15452 ( .A(n7116), .B(n6175), .Z(n6718) );
  HS65_LS_NAND2X2 U15453 ( .A(n5524), .B(n4582), .Z(n5125) );
  HS65_LS_NOR3X1 U15454 ( .A(n1443), .B(n1125), .C(n1387), .Z(n1440) );
  HS65_LS_OAI21X2 U15455 ( .A(n1200), .B(n1173), .C(n1395), .Z(n1443) );
  HS65_LS_NOR3X1 U15456 ( .A(n2195), .B(n1877), .C(n2139), .Z(n2192) );
  HS65_LS_OAI21X2 U15457 ( .A(n1952), .B(n1925), .C(n2147), .Z(n2195) );
  HS65_LS_NOR3X1 U15458 ( .A(n4097), .B(n4098), .C(n3923), .Z(n4094) );
  HS65_LS_OAI21X2 U15459 ( .A(n3057), .B(n3044), .C(n4105), .Z(n4097) );
  HS65_LS_NOR2X2 U15460 ( .A(n3599), .B(n3066), .Z(n3284) );
  HS65_LS_NOR2X2 U15461 ( .A(n2250), .B(n2286), .Z(n2468) );
  HS65_LS_NOR2X2 U15462 ( .A(n1498), .B(n1534), .Z(n1716) );
  HS65_LS_NAND2X2 U15463 ( .A(n45), .B(n4491), .Z(n5059) );
  HS65_LS_NAND2X2 U15464 ( .A(n571), .B(n6084), .Z(n6652) );
  HS65_LS_NAND2X2 U15465 ( .A(n1135), .B(n1153), .Z(n1132) );
  HS65_LS_NAND2X2 U15466 ( .A(n1887), .B(n1905), .Z(n1884) );
  HS65_LS_NAND2X2 U15467 ( .A(n4561), .B(n4559), .Z(n4571) );
  HS65_LS_NAND2X2 U15468 ( .A(n6154), .B(n6152), .Z(n6164) );
  HS65_LS_NOR2X2 U15469 ( .A(n2893), .B(n3173), .Z(n3674) );
  HS65_LS_IVX2 U15470 ( .A(n7761), .Z(n370) );
  HS65_LS_NOR2X2 U15471 ( .A(n1874), .B(n1910), .Z(n2092) );
  HS65_LS_NOR2X2 U15472 ( .A(n1122), .B(n1158), .Z(n1340) );
  HS65_LS_IVX2 U15473 ( .A(n3538), .Z(n193) );
  HS65_LS_NOR2X2 U15474 ( .A(n8040), .B(n7954), .Z(n8516) );
  HS65_LS_IVX2 U15475 ( .A(n1534), .Z(n840) );
  HS65_LS_IVX2 U15476 ( .A(n2286), .Z(n922) );
  HS65_LS_IVX2 U15477 ( .A(n8130), .Z(n387) );
  HS65_LS_NOR2X2 U15478 ( .A(n2842), .B(n3007), .Z(n3873) );
  HS65_LS_NOR2X2 U15479 ( .A(n3726), .B(n3359), .Z(n3781) );
  HS65_LS_NOR2X2 U15480 ( .A(n8571), .B(n8639), .Z(n8383) );
  HS65_LS_NOR2X2 U15481 ( .A(n4002), .B(n3297), .Z(n3659) );
  HS65_LS_NAND2X2 U15482 ( .A(n2855), .B(n3002), .Z(n2852) );
  HS65_LS_NAND2X2 U15483 ( .A(n2900), .B(n2984), .Z(n2897) );
  HS65_LS_NAND2X2 U15484 ( .A(n3905), .B(n3454), .Z(n2872) );
  HS65_LS_IVX2 U15485 ( .A(n2284), .Z(n909) );
  HS65_LS_IVX2 U15486 ( .A(n1156), .Z(n868) );
  HS65_LS_IVX2 U15487 ( .A(n1908), .Z(n786) );
  HS65_LS_IVX2 U15488 ( .A(n1532), .Z(n827) );
  HS65_LS_NAND2X2 U15489 ( .A(n475), .B(n4616), .Z(n5413) );
  HS65_LS_NAND2X2 U15490 ( .A(n298), .B(n6209), .Z(n7005) );
  HS65_LS_NAND2X2 U15491 ( .A(n77), .B(n6184), .Z(n6890) );
  HS65_LS_NAND2X2 U15492 ( .A(n256), .B(n4591), .Z(n5298) );
  HS65_LS_NAND2X2 U15493 ( .A(n527), .B(n6124), .Z(n6773) );
  HS65_LS_NAND2X2 U15494 ( .A(n709), .B(n4531), .Z(n5181) );
  HS65_LS_NOR2X2 U15495 ( .A(n2438), .B(n2342), .Z(n2508) );
  HS65_LS_NOR2X2 U15496 ( .A(n1686), .B(n1590), .Z(n1756) );
  HS65_LS_IVX2 U15497 ( .A(n1910), .Z(n799) );
  HS65_LS_IVX2 U15498 ( .A(n1158), .Z(n881) );
  HS65_LS_NOR2X2 U15499 ( .A(n7857), .B(n7871), .Z(n8289) );
  HS65_LS_IVX2 U15500 ( .A(n3415), .Z(n432) );
  HS65_LS_CBI4I1X3 U15501 ( .A(n2850), .B(n3007), .C(n3415), .D(n3805), .Z(
        n4305) );
  HS65_LS_NAND2X2 U15502 ( .A(n606), .B(n7709), .Z(n8713) );
  HS65_LS_NAND2X2 U15503 ( .A(n119), .B(n7747), .Z(n8801) );
  HS65_LS_NOR2X2 U15504 ( .A(n1310), .B(n1214), .Z(n1380) );
  HS65_LS_NOR2X2 U15505 ( .A(n3148), .B(n3359), .Z(n3160) );
  HS65_LS_NOR2X2 U15506 ( .A(n3189), .B(n3421), .Z(n3201) );
  HS65_LS_IVX2 U15507 ( .A(n7686), .Z(n589) );
  HS65_LS_IVX2 U15508 ( .A(n7724), .Z(n102) );
  HS65_LS_NOR2X2 U15509 ( .A(n8186), .B(n8182), .Z(n7922) );
  HS65_LS_NOR2X2 U15510 ( .A(n8154), .B(n8150), .Z(n7823) );
  HS65_LS_IVX2 U15511 ( .A(n2900), .Z(n646) );
  HS65_LS_IVX2 U15512 ( .A(n3905), .Z(n194) );
  HS65_LS_IVX2 U15513 ( .A(n2855), .Z(n422) );
  HS65_LS_NOR2X2 U15514 ( .A(n2924), .B(n3066), .Z(n3660) );
  HS65_LS_CBI4I1X3 U15515 ( .A(n3415), .B(n3189), .C(n2854), .D(n3830), .Z(
        n3829) );
  HS65_LS_NAND2X2 U15516 ( .A(n133), .B(n7747), .Z(n7901) );
  HS65_LS_NAND2X2 U15517 ( .A(n620), .B(n7709), .Z(n7801) );
  HS65_LS_NAND4ABX3 U15518 ( .A(n8349), .B(n8350), .C(n8351), .D(n8352), .Z(
        n7951) );
  HS65_LS_OAI222X2 U15519 ( .A(n8361), .B(n7960), .C(n8061), .D(n8069), .E(
        n7777), .F(n7779), .Z(n8350) );
  HS65_LS_NOR4ABX2 U15520 ( .A(n8357), .B(n8358), .C(n8359), .D(n8360), .Z(
        n8351) );
  HS65_LS_NAND3X2 U15521 ( .A(n8362), .B(n8363), .C(n8364), .Z(n8349) );
  HS65_LS_NOR2X2 U15522 ( .A(n8639), .B(n7777), .Z(n8620) );
  HS65_LS_NOR2X2 U15523 ( .A(n8663), .B(n7760), .Z(n8231) );
  HS65_LS_NOR2X2 U15524 ( .A(n2062), .B(n1966), .Z(n2132) );
  HS65_LS_IVX2 U15525 ( .A(n8326), .Z(n347) );
  HS65_LS_CBI4I1X3 U15526 ( .A(n8130), .B(n8019), .C(n8252), .D(n8253), .Z(
        n8251) );
  HS65_LS_CBI4I1X3 U15527 ( .A(n8326), .B(n8061), .C(n8556), .D(n8557), .Z(
        n8555) );
  HS65_LS_NAND4ABX3 U15528 ( .A(n8861), .B(n8862), .C(n8863), .D(n8864), .Z(
        n8632) );
  HS65_LS_CBI4I1X3 U15529 ( .A(n7777), .B(n8332), .C(n7961), .D(n8354), .Z(
        n8861) );
  HS65_LS_CBI4I1X3 U15530 ( .A(n355), .B(n8051), .C(n8556), .D(n8873), .Z(
        n8862) );
  HS65_LS_NOR4ABX2 U15531 ( .A(n8617), .B(n8603), .C(n325), .D(n8581), .Z(
        n8863) );
  HS65_LS_IVX2 U15532 ( .A(n2527), .Z(n908) );
  HS65_LS_IVX2 U15533 ( .A(n1775), .Z(n826) );
  HS65_LS_NOR2X2 U15534 ( .A(n3187), .B(n3004), .Z(n3897) );
  HS65_LS_NAND4ABX3 U15535 ( .A(n8652), .B(n8653), .C(n8654), .D(n8655), .Z(
        n8499) );
  HS65_LS_CBI4I1X3 U15536 ( .A(n7760), .B(n8136), .C(n7859), .D(n8112), .Z(
        n8652) );
  HS65_LS_NOR4ABX2 U15537 ( .A(n8234), .B(n8258), .C(n8277), .D(n8300), .Z(
        n8654) );
  HS65_LS_CBI4I1X3 U15538 ( .A(n392), .B(n8009), .C(n8252), .D(n8665), .Z(
        n8653) );
  HS65_LS_NAND2X2 U15539 ( .A(n4784), .B(n4783), .Z(n4794) );
  HS65_LS_NAND2X2 U15540 ( .A(n4745), .B(n4744), .Z(n4755) );
  HS65_LS_NAND2X2 U15541 ( .A(n4638), .B(n4637), .Z(n4648) );
  HS65_LS_NAND2X2 U15542 ( .A(n6377), .B(n6376), .Z(n6387) );
  HS65_LS_NAND2X2 U15543 ( .A(n6338), .B(n6337), .Z(n6348) );
  HS65_LS_NAND2X2 U15544 ( .A(n6231), .B(n6230), .Z(n6241) );
  HS65_LS_NOR2X2 U15545 ( .A(n2986), .B(n3962), .Z(n3170) );
  HS65_LS_NOR2X2 U15546 ( .A(n3484), .B(n3133), .Z(n3542) );
  HS65_LS_NOR2X2 U15547 ( .A(n8018), .B(n7858), .Z(n8318) );
  HS65_LS_NOR2X2 U15548 ( .A(n8060), .B(n7960), .Z(n8534) );
  HS65_LS_NOR2X2 U15549 ( .A(n5041), .B(n4719), .Z(n4727) );
  HS65_LS_NOR2X2 U15550 ( .A(n6634), .B(n6312), .Z(n6320) );
  HS65_LS_NOR2X2 U15551 ( .A(n4669), .B(n4676), .Z(n5127) );
  HS65_LS_NOR2X2 U15552 ( .A(n6262), .B(n6269), .Z(n6720) );
  HS65_LS_NOR2X2 U15553 ( .A(n3297), .B(n3053), .Z(n3645) );
  HS65_LS_NOR2X2 U15554 ( .A(n2989), .B(n3962), .Z(n3356) );
  HS65_LS_NOR2X2 U15555 ( .A(n5395), .B(n4512), .Z(n4995) );
  HS65_LS_NOR2X2 U15556 ( .A(n5280), .B(n4466), .Z(n4941) );
  HS65_LS_NOR2X2 U15557 ( .A(n6987), .B(n6105), .Z(n6588) );
  HS65_LS_NOR2X2 U15558 ( .A(n5163), .B(n4860), .Z(n4867) );
  HS65_LS_NOR2X2 U15559 ( .A(n6755), .B(n6453), .Z(n6460) );
  HS65_LS_NOR2X2 U15560 ( .A(n6872), .B(n6059), .Z(n6534) );
  HS65_LS_NOR2X2 U15561 ( .A(n3281), .B(n3262), .Z(n3285) );
  HS65_LS_OAI21X2 U15562 ( .A(n4680), .B(n4695), .C(n5667), .Z(n5709) );
  HS65_LS_OAI21X2 U15563 ( .A(n6273), .B(n6288), .C(n7259), .Z(n7301) );
  HS65_LS_NAND4ABX3 U15564 ( .A(n9010), .B(n9011), .C(n9012), .D(n9013), .Z(
        n7810) );
  HS65_LS_NOR4ABX2 U15565 ( .A(n8701), .B(n8712), .C(n8758), .D(n8723), .Z(
        n9012) );
  HS65_LS_CB4I6X4 U15566 ( .A(n589), .B(n597), .C(n624), .D(n8415), .Z(n9010)
         );
  HS65_LS_CBI4I1X3 U15567 ( .A(n617), .B(n7633), .C(n7634), .D(n9031), .Z(
        n9011) );
  HS65_LS_NAND4ABX3 U15568 ( .A(n9068), .B(n9069), .C(n9070), .D(n9071), .Z(
        n7910) );
  HS65_LS_NOR4ABX2 U15569 ( .A(n8789), .B(n8800), .C(n8846), .D(n8811), .Z(
        n9070) );
  HS65_LS_CB4I6X4 U15570 ( .A(n102), .B(n110), .C(n137), .D(n8475), .Z(n9068)
         );
  HS65_LS_CBI4I1X3 U15571 ( .A(n130), .B(n7661), .C(n7662), .D(n9089), .Z(
        n9069) );
  HS65_LS_NOR2X2 U15572 ( .A(n1577), .B(n1510), .Z(n1704) );
  HS65_LS_NOR2X2 U15573 ( .A(n2329), .B(n2262), .Z(n2456) );
  HS65_LS_NAND4ABX3 U15574 ( .A(n5557), .B(n5558), .C(n5559), .D(n5560), .Z(
        n4506) );
  HS65_LS_CB4I6X4 U15575 ( .A(n467), .B(n453), .C(n480), .D(n4995), .Z(n5557)
         );
  HS65_LS_NOR4ABX2 U15576 ( .A(n5394), .B(n5412), .C(n5471), .D(n5426), .Z(
        n5559) );
  HS65_LS_CBI4I1X3 U15577 ( .A(n488), .B(n5566), .C(n4516), .D(n5567), .Z(
        n5558) );
  HS65_LS_NAND4ABX3 U15578 ( .A(n5536), .B(n5537), .C(n5538), .D(n5539), .Z(
        n4460) );
  HS65_LS_CB4I6X4 U15579 ( .A(n248), .B(n234), .C(n261), .D(n4941), .Z(n5536)
         );
  HS65_LS_NOR4ABX2 U15580 ( .A(n5279), .B(n5297), .C(n5356), .D(n5311), .Z(
        n5538) );
  HS65_LS_CBI4I1X3 U15581 ( .A(n269), .B(n5545), .C(n4470), .D(n5546), .Z(
        n5537) );
  HS65_LS_NAND4ABX3 U15582 ( .A(n7149), .B(n7150), .C(n7151), .D(n7152), .Z(
        n6099) );
  HS65_LS_CB4I6X4 U15583 ( .A(n290), .B(n276), .C(n303), .D(n6588), .Z(n7149)
         );
  HS65_LS_NOR4ABX2 U15584 ( .A(n6986), .B(n7004), .C(n7063), .D(n7018), .Z(
        n7151) );
  HS65_LS_CBI4I1X3 U15585 ( .A(n311), .B(n7158), .C(n6109), .D(n7159), .Z(
        n7150) );
  HS65_LS_NAND4ABX3 U15586 ( .A(n5789), .B(n5790), .C(n5791), .D(n5792), .Z(
        n5503) );
  HS65_LS_CB4I6X4 U15587 ( .A(n677), .B(n687), .C(n695), .D(n4867), .Z(n5789)
         );
  HS65_LS_NOR4ABX2 U15588 ( .A(n5162), .B(n5180), .C(n5241), .D(n5195), .Z(
        n5791) );
  HS65_LS_CBI4I1X3 U15589 ( .A(n703), .B(n5581), .C(n4535), .D(n5821), .Z(
        n5790) );
  HS65_LS_NAND4ABX3 U15590 ( .A(n5727), .B(n5728), .C(n5729), .D(n5730), .Z(
        n5487) );
  HS65_LS_NOR4ABX2 U15591 ( .A(n5040), .B(n5058), .C(n5105), .D(n5073), .Z(
        n5729) );
  HS65_LS_CBI4I1X3 U15592 ( .A(n39), .B(n5516), .C(n4495), .D(n5759), .Z(n5728) );
  HS65_LS_CB4I6X4 U15593 ( .A(n12), .B(n23), .C(n31), .D(n4727), .Z(n5727) );
  HS65_LS_NAND4ABX3 U15594 ( .A(n7381), .B(n7382), .C(n7383), .D(n7384), .Z(
        n7095) );
  HS65_LS_CB4I6X4 U15595 ( .A(n495), .B(n505), .C(n513), .D(n6460), .Z(n7381)
         );
  HS65_LS_NOR4ABX2 U15596 ( .A(n6754), .B(n6772), .C(n6833), .D(n6787), .Z(
        n7383) );
  HS65_LS_CBI4I1X3 U15597 ( .A(n521), .B(n7173), .C(n6128), .D(n7413), .Z(
        n7382) );
  HS65_LS_NAND4ABX3 U15598 ( .A(n7128), .B(n7129), .C(n7130), .D(n7131), .Z(
        n6053) );
  HS65_LS_CB4I6X4 U15599 ( .A(n69), .B(n55), .C(n82), .D(n6534), .Z(n7128) );
  HS65_LS_NOR4ABX2 U15600 ( .A(n6871), .B(n6889), .C(n6948), .D(n6903), .Z(
        n7130) );
  HS65_LS_CBI4I1X3 U15601 ( .A(n90), .B(n7137), .C(n6063), .D(n7138), .Z(n7129) );
  HS65_LS_NAND4ABX3 U15602 ( .A(n7319), .B(n7320), .C(n7321), .D(n7322), .Z(
        n7079) );
  HS65_LS_NOR4ABX2 U15603 ( .A(n6633), .B(n6651), .C(n6698), .D(n6666), .Z(
        n7321) );
  HS65_LS_CBI4I1X3 U15604 ( .A(n565), .B(n7108), .C(n6088), .D(n7351), .Z(
        n7320) );
  HS65_LS_CB4I6X4 U15605 ( .A(n538), .B(n549), .C(n557), .D(n6320), .Z(n7319)
         );
  HS65_LS_NOR2X2 U15606 ( .A(n8154), .B(n7847), .Z(n8725) );
  HS65_LS_NOR2X2 U15607 ( .A(n8186), .B(n7886), .Z(n8813) );
  HS65_LS_IVX2 U15608 ( .A(n1399), .Z(n867) );
  HS65_LS_NOR2X2 U15609 ( .A(n3146), .B(n2986), .Z(n3780) );
  HS65_LS_OAI21X2 U15610 ( .A(n7760), .B(n8080), .C(n8081), .Z(n8079) );
  HS65_LS_NAND4ABX3 U15611 ( .A(n8107), .B(n8108), .C(n8109), .D(n8110), .Z(
        n7868) );
  HS65_LS_OAI222X2 U15612 ( .A(n8119), .B(n7858), .C(n8019), .D(n8030), .E(
        n7760), .F(n7762), .Z(n8108) );
  HS65_LS_NOR4ABX2 U15613 ( .A(n8111), .B(n8112), .C(n8113), .D(n8114), .Z(
        n8110) );
  HS65_LS_NAND3X2 U15614 ( .A(n8120), .B(n8121), .C(n8122), .Z(n8107) );
  HS65_LS_NOR2X2 U15615 ( .A(n2901), .B(n2989), .Z(n3334) );
  HS65_LS_NOR2X2 U15616 ( .A(n1173), .B(n1214), .Z(n1185) );
  HS65_LS_NOR2X2 U15617 ( .A(n1925), .B(n1966), .Z(n1937) );
  HS65_LS_NOR2X2 U15618 ( .A(n2301), .B(n2342), .Z(n2313) );
  HS65_LS_NOR2X2 U15619 ( .A(n1549), .B(n1590), .Z(n1561) );
  HS65_LS_CBI4I1X3 U15620 ( .A(n7872), .B(n7861), .C(n8130), .D(n8115), .Z(
        n8954) );
  HS65_LS_NOR2X2 U15621 ( .A(n1201), .B(n1134), .Z(n1328) );
  HS65_LS_NOR2X2 U15622 ( .A(n1953), .B(n1886), .Z(n2080) );
  HS65_LS_NOR2X2 U15623 ( .A(n4561), .B(n4676), .Z(n4574) );
  HS65_LS_NOR2X2 U15624 ( .A(n6154), .B(n6269), .Z(n6167) );
  HS65_LS_NOR2X2 U15625 ( .A(n2874), .B(n3940), .Z(n2968) );
  HS65_LS_IVX2 U15626 ( .A(n2151), .Z(n785) );
  HS65_LS_NOR2X2 U15627 ( .A(n5395), .B(n5565), .Z(n5391) );
  HS65_LS_NOR2X2 U15628 ( .A(n5280), .B(n5544), .Z(n5276) );
  HS65_LS_NOR2X2 U15629 ( .A(n5163), .B(n5589), .Z(n5159) );
  HS65_LS_NOR2X2 U15630 ( .A(n6987), .B(n7157), .Z(n6983) );
  HS65_LS_NOR2X2 U15631 ( .A(n6872), .B(n7136), .Z(n6868) );
  HS65_LS_NOR2X2 U15632 ( .A(n6755), .B(n7181), .Z(n6751) );
  HS65_LS_IVX2 U15633 ( .A(n2944), .Z(n217) );
  HS65_LS_IVX2 U15634 ( .A(n3187), .Z(n440) );
  HS65_LS_NOR2X2 U15635 ( .A(n6337), .B(n7210), .Z(n6536) );
  HS65_LS_NOR2X2 U15636 ( .A(n6376), .B(n7237), .Z(n6590) );
  HS65_LS_NOR2X2 U15637 ( .A(n4783), .B(n5645), .Z(n4997) );
  HS65_LS_NOR2X2 U15638 ( .A(n4744), .B(n5618), .Z(n4943) );
  HS65_LS_NOR2X2 U15639 ( .A(n4637), .B(n5591), .Z(n4869) );
  HS65_LS_NOR2X2 U15640 ( .A(n6230), .B(n7183), .Z(n6462) );
  HS65_LS_NOR2X2 U15641 ( .A(n1171), .B(n1155), .Z(n1379) );
  HS65_LS_NOR2X2 U15642 ( .A(n1923), .B(n1907), .Z(n2131) );
  HS65_LS_NOR2X2 U15643 ( .A(n2299), .B(n2283), .Z(n2507) );
  HS65_LS_IVX2 U15644 ( .A(n8149), .Z(n613) );
  HS65_LS_IVX2 U15645 ( .A(n8181), .Z(n126) );
  HS65_LS_NOR2X2 U15646 ( .A(n1547), .B(n1531), .Z(n1755) );
  HS65_LS_NOR2X2 U15647 ( .A(n6059), .B(n6529), .Z(n6499) );
  HS65_LS_NOR2X2 U15648 ( .A(n6105), .B(n6583), .Z(n6553) );
  HS65_LS_NOR2X2 U15649 ( .A(n4466), .B(n4936), .Z(n4906) );
  HS65_LS_NOR2X2 U15650 ( .A(n4512), .B(n4990), .Z(n4960) );
  HS65_LS_NOR2X2 U15651 ( .A(n4860), .B(n4861), .Z(n4829) );
  HS65_LS_NOR2X2 U15652 ( .A(n6453), .B(n6454), .Z(n6422) );
  HS65_LS_NOR2X2 U15653 ( .A(n2946), .B(n3133), .Z(n2957) );
  HS65_LS_CBI4I1X3 U15654 ( .A(n7955), .B(n7963), .C(n8326), .D(n8357), .Z(
        n8894) );
  HS65_LS_OAI21X2 U15655 ( .A(n7777), .B(n8335), .C(n8336), .Z(n8334) );
  HS65_LS_IVX2 U15656 ( .A(n8379), .Z(n354) );
  HS65_LS_NOR2X2 U15657 ( .A(n7778), .B(n8051), .Z(n8625) );
  HS65_LS_NOR2X2 U15658 ( .A(n2944), .B(n2874), .Z(n3540) );
  HS65_LS_NOR2X2 U15659 ( .A(n3209), .B(n2854), .Z(n3861) );
  HS65_LS_IVX2 U15660 ( .A(n8315), .Z(n395) );
  HS65_LS_IVX2 U15661 ( .A(n3486), .Z(n205) );
  HS65_LS_IVX2 U15662 ( .A(n7961), .Z(n345) );
  HS65_LS_NAND4ABX3 U15663 ( .A(n2381), .B(n2382), .C(n2383), .D(n2384), .Z(
        n2277) );
  HS65_LS_NOR3X1 U15664 ( .A(n2385), .B(n2386), .C(n2387), .Z(n2384) );
  HS65_LS_AOI222X2 U15665 ( .A(n920), .B(n900), .C(n918), .D(n901), .E(n924), 
        .F(n905), .Z(n2383) );
  HS65_LS_OAI212X3 U15666 ( .A(n2391), .B(n2250), .C(n2323), .D(n2264), .E(
        n2392), .Z(n2381) );
  HS65_LS_NAND4ABX3 U15667 ( .A(n1629), .B(n1630), .C(n1631), .D(n1632), .Z(
        n1525) );
  HS65_LS_NOR3X1 U15668 ( .A(n1633), .B(n1634), .C(n1635), .Z(n1632) );
  HS65_LS_AOI222X2 U15669 ( .A(n838), .B(n818), .C(n836), .D(n819), .E(n842), 
        .F(n823), .Z(n1631) );
  HS65_LS_OAI212X3 U15670 ( .A(n1639), .B(n1498), .C(n1571), .D(n1512), .E(
        n1640), .Z(n1629) );
  HS65_LS_NOR2X2 U15671 ( .A(n6059), .B(n6051), .Z(n6349) );
  HS65_LS_NOR2X2 U15672 ( .A(n4512), .B(n4504), .Z(n4795) );
  HS65_LS_NOR2X2 U15673 ( .A(n6105), .B(n6097), .Z(n6388) );
  HS65_LS_NOR2X2 U15674 ( .A(n4466), .B(n4458), .Z(n4756) );
  HS65_LS_NOR2X2 U15675 ( .A(n4860), .B(n4820), .Z(n4649) );
  HS65_LS_NOR2X2 U15676 ( .A(n6453), .B(n6413), .Z(n6242) );
  HS65_LS_NAND4ABX3 U15677 ( .A(n1253), .B(n1254), .C(n1255), .D(n1256), .Z(
        n1149) );
  HS65_LS_NOR3X1 U15678 ( .A(n1257), .B(n1258), .C(n1259), .Z(n1256) );
  HS65_LS_AOI222X2 U15679 ( .A(n879), .B(n859), .C(n877), .D(n860), .E(n883), 
        .F(n864), .Z(n1255) );
  HS65_LS_OAI212X3 U15680 ( .A(n1263), .B(n1122), .C(n1195), .D(n1136), .E(
        n1264), .Z(n1253) );
  HS65_LS_NAND4ABX3 U15681 ( .A(n2005), .B(n2006), .C(n2007), .D(n2008), .Z(
        n1901) );
  HS65_LS_NOR3X1 U15682 ( .A(n2009), .B(n2010), .C(n2011), .Z(n2008) );
  HS65_LS_AOI222X2 U15683 ( .A(n797), .B(n777), .C(n795), .D(n778), .E(n801), 
        .F(n782), .Z(n2007) );
  HS65_LS_OAI212X3 U15684 ( .A(n2015), .B(n1874), .C(n1947), .D(n1888), .E(
        n2016), .Z(n2005) );
  HS65_LS_NAND2X2 U15685 ( .A(n3845), .B(n3004), .Z(n3787) );
  HS65_LS_NOR2X2 U15686 ( .A(n5041), .B(n5524), .Z(n5037) );
  HS65_LS_NOR2X2 U15687 ( .A(n6634), .B(n7116), .Z(n6630) );
  HS65_LS_AOI12X2 U15688 ( .A(n2841), .B(n3845), .C(n3843), .Z(n3984) );
  HS65_LS_NOR2X2 U15689 ( .A(n3052), .B(n3262), .Z(n3655) );
  HS65_LS_NOR2X2 U15690 ( .A(n7842), .B(n8699), .Z(n8415) );
  HS65_LS_NOR2X2 U15691 ( .A(n7881), .B(n8787), .Z(n8475) );
  HS65_LS_NOR2X2 U15692 ( .A(n7959), .B(n8639), .Z(n8573) );
  HS65_LS_IVX2 U15693 ( .A(n7872), .Z(n366) );
  HS65_LS_NOR2X2 U15694 ( .A(n3263), .B(n3262), .Z(n3287) );
  HS65_LS_NAND2X2 U15695 ( .A(n8267), .B(n7858), .Z(n8208) );
  HS65_LS_NAND2X2 U15696 ( .A(n8571), .B(n7960), .Z(n8513) );
  HS65_LS_NOR2X2 U15697 ( .A(n7861), .B(n8119), .Z(n8283) );
  HS65_LS_IVX2 U15698 ( .A(n7670), .Z(n98) );
  HS65_LS_IVX2 U15699 ( .A(n7642), .Z(n585) );
  HS65_LS_NAND2X2 U15700 ( .A(n3728), .B(n2986), .Z(n3670) );
  HS65_LS_NOR2X2 U15701 ( .A(n3843), .B(n3421), .Z(n3898) );
  HS65_LS_NOR2X2 U15702 ( .A(n4577), .B(n4721), .Z(n5102) );
  HS65_LS_NOR2X2 U15703 ( .A(n6170), .B(n6314), .Z(n6695) );
  HS65_LS_NOR2X2 U15704 ( .A(n4784), .B(n5008), .Z(n4797) );
  HS65_LS_NOR2X2 U15705 ( .A(n4745), .B(n4894), .Z(n4758) );
  HS65_LS_NOR2X2 U15706 ( .A(n6377), .B(n6601), .Z(n6390) );
  HS65_LS_NOR2X2 U15707 ( .A(n6338), .B(n6487), .Z(n6351) );
  HS65_LS_NOR2X2 U15708 ( .A(n4638), .B(n4880), .Z(n4651) );
  HS65_LS_NOR2X2 U15709 ( .A(n6231), .B(n6473), .Z(n6244) );
  HS65_LS_NOR2X2 U15710 ( .A(n3168), .B(n2899), .Z(n3744) );
  HS65_LS_NOR2X2 U15711 ( .A(n3065), .B(n3057), .Z(n3621) );
  HS65_LS_IVX2 U15712 ( .A(n2887), .Z(n669) );
  HS65_LS_IVX2 U15713 ( .A(n3281), .Z(n148) );
  HS65_LS_NOR2X2 U15714 ( .A(n2848), .B(n3415), .Z(n3789) );
  HS65_LS_IVX2 U15715 ( .A(n3066), .Z(n171) );
  HS65_LS_OAI21X2 U15716 ( .A(n3421), .B(n2849), .C(n3796), .Z(n4321) );
  HS65_LS_NOR2X2 U15717 ( .A(n8159), .B(n7842), .Z(n8424) );
  HS65_LS_NOR2X2 U15718 ( .A(n8191), .B(n7881), .Z(n8484) );
  HS65_LS_NOR2X2 U15719 ( .A(n7697), .B(n7633), .Z(n8165) );
  HS65_LS_NOR2X2 U15720 ( .A(n7735), .B(n7661), .Z(n8197) );
  HS65_LS_IVX2 U15721 ( .A(n7870), .Z(n372) );
  HS65_LS_NAND2X2 U15722 ( .A(n8671), .B(n7859), .Z(n8506) );
  HS65_LS_IVX2 U15723 ( .A(n8267), .Z(n375) );
  HS65_LS_NAND2X2 U15724 ( .A(n1312), .B(n1155), .Z(n1270) );
  HS65_LS_NAND2X2 U15725 ( .A(n2064), .B(n1907), .Z(n2022) );
  HS65_LS_NAND2X2 U15726 ( .A(n2440), .B(n2283), .Z(n2398) );
  HS65_LS_NOR2X2 U15727 ( .A(n2925), .B(n3057), .Z(n3654) );
  HS65_LS_NOR2X2 U15728 ( .A(n8267), .B(n8663), .Z(n8089) );
  HS65_LS_NAND2X2 U15729 ( .A(n1688), .B(n1531), .Z(n1646) );
  HS65_LS_NOR2X2 U15730 ( .A(n6273), .B(n6312), .Z(n6165) );
  HS65_LS_NOR2X2 U15731 ( .A(n4680), .B(n4719), .Z(n4572) );
  HS65_LS_IVX2 U15732 ( .A(n3146), .Z(n664) );
  HS65_LS_NOR2X2 U15733 ( .A(n5002), .B(n5008), .Z(n4520) );
  HS65_LS_NOR2X2 U15734 ( .A(n4888), .B(n4894), .Z(n4474) );
  HS65_LS_NOR2X2 U15735 ( .A(n6595), .B(n6601), .Z(n6113) );
  HS65_LS_NOR2X2 U15736 ( .A(n4874), .B(n4880), .Z(n5233) );
  HS65_LS_NOR2X2 U15737 ( .A(n6467), .B(n6473), .Z(n6825) );
  HS65_LS_NOR2X2 U15738 ( .A(n6481), .B(n6487), .Z(n6067) );
  HS65_LS_NOR4ABX2 U15739 ( .A(n7076), .B(n7105), .C(n7106), .D(n7107), .Z(
        n7104) );
  HS65_LS_OAI212X3 U15740 ( .A(n7108), .B(n6153), .C(n7109), .D(n6088), .E(
        n7110), .Z(n7107) );
  HS65_LS_NOR4ABX2 U15741 ( .A(n5484), .B(n5513), .C(n5514), .D(n5515), .Z(
        n5512) );
  HS65_LS_OAI212X3 U15742 ( .A(n5516), .B(n4560), .C(n5517), .D(n4495), .E(
        n5518), .Z(n5515) );
  HS65_LS_IVX2 U15743 ( .A(n2877), .Z(n204) );
  HS65_LS_IVX2 U15744 ( .A(n2989), .Z(n636) );
  HS65_LS_NOR2X2 U15745 ( .A(n4719), .B(n4721), .Z(n4688) );
  HS65_LS_NOR2X2 U15746 ( .A(n6312), .B(n6314), .Z(n6281) );
  HS65_LS_NOR2X2 U15747 ( .A(n7857), .B(n8119), .Z(n8027) );
  HS65_LS_NOR2X2 U15748 ( .A(n7817), .B(n7638), .Z(n8682) );
  HS65_LS_NOR2X2 U15749 ( .A(n7880), .B(n7666), .Z(n8770) );
  HS65_LS_IVX2 U15750 ( .A(n5524), .Z(n48) );
  HS65_LS_IVX2 U15751 ( .A(n7116), .Z(n574) );
  HS65_LS_IVX2 U15752 ( .A(n5565), .Z(n472) );
  HS65_LS_IVX2 U15753 ( .A(n7157), .Z(n295) );
  HS65_LS_IVX2 U15754 ( .A(n7136), .Z(n74) );
  HS65_LS_IVX2 U15755 ( .A(n5544), .Z(n253) );
  HS65_LS_IVX2 U15756 ( .A(n5589), .Z(n712) );
  HS65_LS_IVX2 U15757 ( .A(n7181), .Z(n530) );
  HS65_LS_NOR4ABX2 U15758 ( .A(n3142), .B(n3143), .C(n3144), .D(n3145), .Z(
        n2978) );
  HS65_LS_OAI212X3 U15759 ( .A(n2895), .B(n3146), .C(n3147), .D(n3148), .E(
        n3149), .Z(n3145) );
  HS65_LS_NAND3AX3 U15760 ( .A(n3150), .B(n3151), .C(n3152), .Z(n3144) );
  HS65_LS_NOR3AX2 U15761 ( .A(n3158), .B(n3159), .C(n3160), .Z(n3142) );
  HS65_LS_IVX2 U15762 ( .A(n8332), .Z(n331) );
  HS65_LS_NAND2X2 U15763 ( .A(n3486), .B(n2874), .Z(n3426) );
  HS65_LS_IVX2 U15764 ( .A(n7846), .Z(n584) );
  HS65_LS_IVX2 U15765 ( .A(n7885), .Z(n97) );
  HS65_LS_IVX2 U15766 ( .A(n8119), .Z(n397) );
  HS65_LS_NOR4ABX2 U15767 ( .A(n3274), .B(n3275), .C(n3276), .D(n3277), .Z(
        n2916) );
  HS65_LS_OAI222X2 U15768 ( .A(n3280), .B(n3281), .C(n3282), .D(n3264), .E(
        n3057), .F(n3053), .Z(n3276) );
  HS65_LS_OAI212X3 U15769 ( .A(n3278), .B(n3064), .C(n3236), .D(n3052), .E(
        n3279), .Z(n3277) );
  HS65_LS_NOR3AX2 U15770 ( .A(n3283), .B(n3284), .C(n3285), .Z(n3275) );
  HS65_LS_IVX2 U15771 ( .A(n3893), .Z(n447) );
  HS65_LS_IVX2 U15772 ( .A(n1547), .Z(n825) );
  HS65_LS_IVX2 U15773 ( .A(n2299), .Z(n907) );
  HS65_LS_NOR2X2 U15774 ( .A(n2842), .B(n3845), .Z(n3860) );
  HS65_LS_OAI21X2 U15775 ( .A(n8119), .B(n8136), .C(n8233), .Z(n8960) );
  HS65_LS_NOR2X2 U15776 ( .A(n7645), .B(n8699), .Z(n8426) );
  HS65_LS_NOR2X2 U15777 ( .A(n7673), .B(n8787), .Z(n8486) );
  HS65_LS_NAND2X2 U15778 ( .A(n6634), .B(n6313), .Z(n6607) );
  HS65_LS_NAND2X2 U15779 ( .A(n5041), .B(n4720), .Z(n5014) );
  HS65_LS_NAND2X2 U15780 ( .A(n6872), .B(n6528), .Z(n6846) );
  HS65_LS_NAND2X2 U15781 ( .A(n5280), .B(n4935), .Z(n5254) );
  HS65_LS_NAND2X2 U15782 ( .A(n5395), .B(n4989), .Z(n5369) );
  HS65_LS_NAND2X2 U15783 ( .A(n6987), .B(n6582), .Z(n6961) );
  HS65_LS_NAND2X2 U15784 ( .A(n6755), .B(n6452), .Z(n6728) );
  HS65_LS_NAND2X2 U15785 ( .A(n5163), .B(n4859), .Z(n5136) );
  HS65_LS_NOR2X2 U15786 ( .A(n2928), .B(n3058), .Z(n3569) );
  HS65_LS_NOR4ABX2 U15787 ( .A(n3183), .B(n3184), .C(n3185), .D(n3186), .Z(
        n2996) );
  HS65_LS_OAI212X3 U15788 ( .A(n2850), .B(n3187), .C(n3188), .D(n3189), .E(
        n3190), .Z(n3186) );
  HS65_LS_NAND3AX3 U15789 ( .A(n3191), .B(n3192), .C(n3193), .Z(n3185) );
  HS65_LS_NOR4ABX2 U15790 ( .A(n3195), .B(n3196), .C(n3197), .D(n3198), .Z(
        n3184) );
  HS65_LS_IVX2 U15791 ( .A(n7191), .Z(n87) );
  HS65_LS_IVX2 U15792 ( .A(n5599), .Z(n266) );
  HS65_LS_IVX2 U15793 ( .A(n5626), .Z(n485) );
  HS65_LS_IVX2 U15794 ( .A(n7218), .Z(n308) );
  HS65_LS_IVX2 U15795 ( .A(n7174), .Z(n525) );
  HS65_LS_IVX2 U15796 ( .A(n5582), .Z(n707) );
  HS65_LS_OAI21X2 U15797 ( .A(n3359), .B(n2894), .C(n3679), .Z(n4262) );
  HS65_LS_NOR4ABX2 U15798 ( .A(n2939), .B(n2940), .C(n2941), .D(n2942), .Z(
        n2866) );
  HS65_LS_OAI212X3 U15799 ( .A(n2943), .B(n2944), .C(n2945), .D(n2946), .E(
        n2947), .Z(n2942) );
  HS65_LS_NAND3AX3 U15800 ( .A(n2948), .B(n2949), .C(n2950), .Z(n2941) );
  HS65_LS_NOR3AX2 U15801 ( .A(n2956), .B(n2957), .C(n2958), .Z(n2939) );
  HS65_LS_OAI21X2 U15802 ( .A(n3133), .B(n3100), .C(n3435), .Z(n4218) );
  HS65_LS_NOR2X2 U15803 ( .A(n1775), .B(n1571), .Z(n1649) );
  HS65_LS_NOR2X2 U15804 ( .A(n2527), .B(n2323), .Z(n2401) );
  HS65_LS_IVX2 U15805 ( .A(n3123), .Z(n223) );
  HS65_LS_NAND3X2 U15806 ( .A(n1775), .B(n1584), .C(n1570), .Z(n1805) );
  HS65_LS_NAND3X2 U15807 ( .A(n2527), .B(n2336), .C(n2322), .Z(n2557) );
  HS65_LS_NOR2X2 U15808 ( .A(n2314), .B(n2250), .Z(n2312) );
  HS65_LS_NOR2X2 U15809 ( .A(n1562), .B(n1498), .Z(n1560) );
  HS65_LS_NOR2X2 U15810 ( .A(n3282), .B(n3053), .Z(n3622) );
  HS65_LS_IVX2 U15811 ( .A(n1171), .Z(n866) );
  HS65_LS_IVX2 U15812 ( .A(n4835), .Z(n706) );
  HS65_LS_IVX2 U15813 ( .A(n4503), .Z(n489) );
  HS65_LS_IVX2 U15814 ( .A(n6096), .Z(n312) );
  HS65_LS_IVX2 U15815 ( .A(n6050), .Z(n91) );
  HS65_LS_IVX2 U15816 ( .A(n6428), .Z(n524) );
  HS65_LS_IVX2 U15817 ( .A(n4457), .Z(n270) );
  HS65_LS_IVX2 U15818 ( .A(n3262), .Z(n169) );
  HS65_LS_IVX2 U15819 ( .A(n2849), .Z(n442) );
  HS65_LS_NAND3X2 U15820 ( .A(n1399), .B(n1208), .C(n1194), .Z(n1429) );
  HS65_LS_NAND3X2 U15821 ( .A(n2151), .B(n1960), .C(n1946), .Z(n2181) );
  HS65_LS_NOR2X2 U15822 ( .A(n1122), .B(n1312), .Z(n1327) );
  HS65_LS_NOR2X2 U15823 ( .A(n1874), .B(n2064), .Z(n2079) );
  HS65_LS_NOR2X2 U15824 ( .A(n1186), .B(n1122), .Z(n1184) );
  HS65_LS_NOR2X2 U15825 ( .A(n1938), .B(n1874), .Z(n1936) );
  HS65_LS_NOR4ABX2 U15826 ( .A(n3949), .B(n4010), .C(n2891), .D(n4011), .Z(
        n4009) );
  HS65_LS_OA212X4 U15827 ( .A(n2895), .B(n3174), .C(n3776), .D(n2899), .E(
        n3959), .Z(n4010) );
  HS65_LS_NOR2X2 U15828 ( .A(n1498), .B(n1688), .Z(n1703) );
  HS65_LS_NOR2X2 U15829 ( .A(n2250), .B(n2440), .Z(n2455) );
  HS65_LS_NOR4ABX2 U15830 ( .A(n7628), .B(n7629), .C(n7630), .D(n7631), .Z(
        n7627) );
  HS65_LS_OA212X4 U15831 ( .A(n7632), .B(n7633), .C(n7634), .D(n7635), .E(
        n7636), .Z(n7629) );
  HS65_LS_NOR4ABX2 U15832 ( .A(n7656), .B(n7657), .C(n7658), .D(n7659), .Z(
        n7655) );
  HS65_LS_OA212X4 U15833 ( .A(n7660), .B(n7661), .C(n7662), .D(n7663), .E(
        n7664), .Z(n7657) );
  HS65_LS_NOR4ABX2 U15834 ( .A(n3970), .B(n4034), .C(n2846), .D(n4035), .Z(
        n4033) );
  HS65_LS_OA212X4 U15835 ( .A(n2850), .B(n3215), .C(n3893), .D(n2854), .E(
        n3980), .Z(n4034) );
  HS65_LS_NOR2X2 U15836 ( .A(n2151), .B(n1947), .Z(n2025) );
  HS65_LS_NOR2X2 U15837 ( .A(n1399), .B(n1195), .Z(n1273) );
  HS65_LS_IVX2 U15838 ( .A(n7666), .Z(n122) );
  HS65_LS_IVX2 U15839 ( .A(n7638), .Z(n609) );
  HS65_LS_NOR2X2 U15840 ( .A(n3123), .B(n3486), .Z(n3502) );
  HS65_LS_IVX2 U15841 ( .A(n7955), .Z(n321) );
  HS65_LS_IVX2 U15842 ( .A(n1923), .Z(n784) );
  HS65_LS_NOR2X2 U15843 ( .A(n2282), .B(n2250), .Z(n2385) );
  HS65_LS_NOR2X2 U15844 ( .A(n1530), .B(n1498), .Z(n1633) );
  HS65_LS_NAND2X2 U15845 ( .A(n7136), .B(n6359), .Z(n6939) );
  HS65_LS_NAND2X2 U15846 ( .A(n5544), .B(n4766), .Z(n5347) );
  HS65_LS_NAND2X2 U15847 ( .A(n5565), .B(n4805), .Z(n5462) );
  HS65_LS_NAND2X2 U15848 ( .A(n7157), .B(n6398), .Z(n7054) );
  HS65_LS_NAND2X2 U15849 ( .A(n7181), .B(n6252), .Z(n6823) );
  HS65_LS_NAND2X2 U15850 ( .A(n5589), .B(n4659), .Z(n5231) );
  HS65_LS_IVX2 U15851 ( .A(n1214), .Z(n875) );
  HS65_LS_IVX2 U15852 ( .A(n1966), .Z(n793) );
  HS65_LS_IVX2 U15853 ( .A(n2342), .Z(n916) );
  HS65_LS_IVX2 U15854 ( .A(n1590), .Z(n834) );
  HS65_LS_NOR2X2 U15855 ( .A(n8332), .B(n8061), .Z(n8073) );
  HS65_LS_IVX2 U15856 ( .A(n6312), .Z(n561) );
  HS65_LS_IVX2 U15857 ( .A(n4719), .Z(n35) );
  HS65_LS_NOR2X2 U15858 ( .A(n3538), .B(n3123), .Z(n2958) );
  HS65_LS_IVX2 U15859 ( .A(n6059), .Z(n86) );
  HS65_LS_IVX2 U15860 ( .A(n4512), .Z(n484) );
  HS65_LS_IVX2 U15861 ( .A(n6105), .Z(n307) );
  HS65_LS_IVX2 U15862 ( .A(n4466), .Z(n265) );
  HS65_LS_IVX2 U15863 ( .A(n4860), .Z(n699) );
  HS65_LS_IVX2 U15864 ( .A(n6453), .Z(n517) );
  HS65_LS_NOR2X2 U15865 ( .A(n2887), .B(n3728), .Z(n3743) );
  HS65_LS_NOR2X2 U15866 ( .A(n1584), .B(n1590), .Z(n1514) );
  HS65_LS_NOR2X2 U15867 ( .A(n2336), .B(n2342), .Z(n2266) );
  HS65_LS_IVX2 U15868 ( .A(n7632), .Z(n592) );
  HS65_LS_IVX2 U15869 ( .A(n7660), .Z(n105) );
  HS65_LS_IVX2 U15870 ( .A(n3776), .Z(n671) );
  HS65_LS_NOR2X2 U15871 ( .A(n1154), .B(n1122), .Z(n1257) );
  HS65_LS_NOR2X2 U15872 ( .A(n1906), .B(n1874), .Z(n2009) );
  HS65_LS_IVX2 U15873 ( .A(n4783), .Z(n482) );
  HS65_LS_IVX2 U15874 ( .A(n4744), .Z(n263) );
  HS65_LS_IVX2 U15875 ( .A(n4637), .Z(n702) );
  HS65_LS_IVX2 U15876 ( .A(n6376), .Z(n305) );
  HS65_LS_IVX2 U15877 ( .A(n6337), .Z(n84) );
  HS65_LS_IVX2 U15878 ( .A(n6230), .Z(n520) );
  HS65_LS_NAND3X2 U15879 ( .A(n3173), .B(n3353), .C(n3161), .Z(n4028) );
  HS65_LS_NOR2X2 U15880 ( .A(n1208), .B(n1214), .Z(n1138) );
  HS65_LS_NOR2X2 U15881 ( .A(n7778), .B(n8379), .Z(n8072) );
  HS65_LS_IVX2 U15882 ( .A(n4559), .Z(n38) );
  HS65_LS_IVX2 U15883 ( .A(n6152), .Z(n564) );
  HS65_LS_NOR2X2 U15884 ( .A(n3778), .B(n2887), .Z(n3159) );
  HS65_LS_NAND2X2 U15885 ( .A(n8881), .B(n7961), .Z(n8644) );
  HS65_LS_NOR2X2 U15886 ( .A(n8070), .B(n8556), .Z(n8527) );
  HS65_LS_NAND2X2 U15887 ( .A(n7686), .B(n7697), .Z(n7684) );
  HS65_LS_NAND2X2 U15888 ( .A(n7724), .B(n7735), .Z(n7722) );
  HS65_LS_NOR2X2 U15889 ( .A(n2873), .B(n3123), .Z(n3116) );
  HS65_LS_NOR2X2 U15890 ( .A(n1960), .B(n1966), .Z(n1890) );
  HS65_LS_NOR2X2 U15891 ( .A(n5395), .B(n4783), .Z(n5397) );
  HS65_LS_NOR2X2 U15892 ( .A(n5280), .B(n4744), .Z(n5282) );
  HS65_LS_NOR2X2 U15893 ( .A(n6987), .B(n6376), .Z(n6989) );
  HS65_LS_NOR2X2 U15894 ( .A(n5163), .B(n4637), .Z(n5165) );
  HS65_LS_NOR2X2 U15895 ( .A(n6755), .B(n6230), .Z(n6757) );
  HS65_LS_NOR2X2 U15896 ( .A(n6872), .B(n6337), .Z(n6874) );
  HS65_LS_NOR4ABX2 U15897 ( .A(n8014), .B(n8015), .C(n8016), .D(n8017), .Z(
        n7866) );
  HS65_LS_OAI212X3 U15898 ( .A(n8018), .B(n7872), .C(n8019), .D(n8004), .E(
        n8020), .Z(n8017) );
  HS65_LS_NOR3X1 U15899 ( .A(n7757), .B(n8028), .C(n8029), .Z(n8014) );
  HS65_LS_NAND4ABX3 U15900 ( .A(n8021), .B(n8022), .C(n8023), .D(n8024), .Z(
        n8016) );
  HS65_LS_NAND3X2 U15901 ( .A(n7638), .B(n7639), .C(n7640), .Z(n7637) );
  HS65_LS_NAND3X2 U15902 ( .A(n7666), .B(n7667), .C(n7668), .Z(n7665) );
  HS65_LS_NAND2X2 U15903 ( .A(n7778), .B(n7953), .Z(n8522) );
  HS65_LS_NOR2X2 U15904 ( .A(n3353), .B(n3359), .Z(n2903) );
  HS65_LS_NOR4ABX2 U15905 ( .A(n8656), .B(n8497), .C(n8651), .D(n8948), .Z(
        n8947) );
  HS65_LS_OAI212X3 U15906 ( .A(n8009), .B(n7872), .C(n8252), .D(n8315), .E(
        n7764), .Z(n8948) );
  HS65_LS_IVX2 U15907 ( .A(n7778), .Z(n335) );
  HS65_LS_NAND2X2 U15908 ( .A(n3281), .B(n3282), .Z(n3596) );
  HS65_LS_NOR2X2 U15909 ( .A(n5041), .B(n4559), .Z(n5043) );
  HS65_LS_NOR2X2 U15910 ( .A(n6634), .B(n6152), .Z(n6636) );
  HS65_LS_NOR2X2 U15911 ( .A(n6354), .B(n6529), .Z(n6945) );
  HS65_LS_NOR2X2 U15912 ( .A(n6247), .B(n6454), .Z(n6830) );
  HS65_LS_NOR2X2 U15913 ( .A(n4654), .B(n4861), .Z(n5238) );
  HS65_LS_NOR2X2 U15914 ( .A(n4800), .B(n4990), .Z(n5468) );
  HS65_LS_NOR2X2 U15915 ( .A(n6393), .B(n6583), .Z(n7060) );
  HS65_LS_NOR2X2 U15916 ( .A(n4761), .B(n4936), .Z(n5353) );
  HS65_LS_IVX2 U15917 ( .A(n2850), .Z(n426) );
  HS65_LS_IVX2 U15918 ( .A(n2894), .Z(n666) );
  HS65_LS_IVX2 U15919 ( .A(n3100), .Z(n215) );
  HS65_LS_AOI12X2 U15920 ( .A(n6194), .B(n6487), .C(n6488), .Z(n6483) );
  HS65_LS_AOI12X2 U15921 ( .A(n6206), .B(n6601), .C(n6602), .Z(n6597) );
  HS65_LS_AOI12X2 U15922 ( .A(n4601), .B(n4894), .C(n4895), .Z(n4890) );
  HS65_LS_AOI12X2 U15923 ( .A(n4613), .B(n5008), .C(n5009), .Z(n5004) );
  HS65_LS_NOR2X2 U15924 ( .A(n7857), .B(n8663), .Z(n8269) );
  HS65_LS_NAND4ABX3 U15925 ( .A(n8392), .B(n8393), .C(n8394), .D(n8395), .Z(
        n8144) );
  HS65_LS_NAND4ABX3 U15926 ( .A(n7798), .B(n8416), .C(n8417), .D(n8418), .Z(
        n8393) );
  HS65_LS_NOR4ABX2 U15927 ( .A(n8396), .B(n8397), .C(n8398), .D(n8399), .Z(
        n8395) );
  HS65_LS_MX41X4 U15928 ( .D0(n614), .S0(n7709), .D1(n592), .S1(n620), .D2(
        n606), .S2(n600), .D3(n594), .S3(n616), .Z(n8392) );
  HS65_LS_NAND4ABX3 U15929 ( .A(n8452), .B(n8453), .C(n8454), .D(n8455), .Z(
        n8176) );
  HS65_LS_NAND4ABX3 U15930 ( .A(n7898), .B(n8476), .C(n8477), .D(n8478), .Z(
        n8453) );
  HS65_LS_NOR4ABX2 U15931 ( .A(n8456), .B(n8457), .C(n8458), .D(n8459), .Z(
        n8455) );
  HS65_LS_MX41X4 U15932 ( .D0(n127), .S0(n7747), .D1(n105), .S1(n133), .D2(
        n119), .S2(n113), .D3(n107), .S3(n129), .Z(n8452) );
  HS65_LS_NOR4ABX2 U15933 ( .A(n7125), .B(n7133), .C(n6055), .D(n7190), .Z(
        n7189) );
  HS65_LS_OAI212X3 U15934 ( .A(n7137), .B(n6058), .C(n7191), .D(n6063), .E(
        n7192), .Z(n7190) );
  HS65_LS_NOR4ABX2 U15935 ( .A(n5554), .B(n5562), .C(n4508), .D(n5625), .Z(
        n5624) );
  HS65_LS_OAI212X3 U15936 ( .A(n5566), .B(n4511), .C(n5626), .D(n4516), .E(
        n5627), .Z(n5625) );
  HS65_LS_NOR4ABX2 U15937 ( .A(n7146), .B(n7154), .C(n6101), .D(n7217), .Z(
        n7216) );
  HS65_LS_OAI212X3 U15938 ( .A(n7158), .B(n6104), .C(n7218), .D(n6109), .E(
        n7219), .Z(n7217) );
  HS65_LS_NOR4ABX2 U15939 ( .A(n5533), .B(n5541), .C(n4462), .D(n5598), .Z(
        n5597) );
  HS65_LS_OAI212X3 U15940 ( .A(n5545), .B(n4465), .C(n5599), .D(n4470), .E(
        n5600), .Z(n5598) );
  HS65_LS_NOR4ABX2 U15941 ( .A(n5500), .B(n5578), .C(n5579), .D(n5580), .Z(
        n5577) );
  HS65_LS_OAI212X3 U15942 ( .A(n5581), .B(n4636), .C(n5582), .D(n4535), .E(
        n5583), .Z(n5580) );
  HS65_LS_NOR4ABX2 U15943 ( .A(n7092), .B(n7170), .C(n7171), .D(n7172), .Z(
        n7169) );
  HS65_LS_OAI212X3 U15944 ( .A(n7173), .B(n6229), .C(n7174), .D(n6128), .E(
        n7175), .Z(n7172) );
  HS65_LS_NOR4ABX2 U15945 ( .A(n8056), .B(n8057), .C(n8058), .D(n8059), .Z(
        n7949) );
  HS65_LS_OAI212X3 U15946 ( .A(n8060), .B(n7955), .C(n8061), .D(n8046), .E(
        n8062), .Z(n8059) );
  HS65_LS_NOR3X1 U15947 ( .A(n8071), .B(n8072), .C(n8073), .Z(n8056) );
  HS65_LS_NAND4ABX3 U15948 ( .A(n8063), .B(n8064), .C(n8065), .D(n8066), .Z(
        n8058) );
  HS65_LS_NOR2X2 U15949 ( .A(n3003), .B(n2842), .Z(n3405) );
  HS65_LS_NOR2X2 U15950 ( .A(n7662), .B(n7932), .Z(n8825) );
  HS65_LS_NOR2X2 U15951 ( .A(n7634), .B(n7833), .Z(n8737) );
  HS65_LS_NOR2X2 U15952 ( .A(n3101), .B(n2971), .Z(n2948) );
  HS65_LS_NAND4ABX3 U15953 ( .A(n6506), .B(n6507), .C(n6508), .D(n6509), .Z(
        n6332) );
  HS65_LS_NAND4ABX3 U15954 ( .A(n6535), .B(n6536), .C(n6537), .D(n6538), .Z(
        n6507) );
  HS65_LS_NOR4ABX2 U15955 ( .A(n6510), .B(n6511), .C(n6512), .D(n6513), .Z(
        n6509) );
  HS65_LS_MX41X4 U15956 ( .D0(n6184), .S0(n85), .D1(n70), .S1(n87), .D2(n77), 
        .S2(n59), .D3(n56), .S3(n89), .Z(n6506) );
  HS65_LS_NAND4ABX3 U15957 ( .A(n6560), .B(n6561), .C(n6562), .D(n6563), .Z(
        n6371) );
  HS65_LS_NAND4ABX3 U15958 ( .A(n6589), .B(n6590), .C(n6591), .D(n6592), .Z(
        n6561) );
  HS65_LS_NOR4ABX2 U15959 ( .A(n6564), .B(n6565), .C(n6566), .D(n6567), .Z(
        n6563) );
  HS65_LS_MX41X4 U15960 ( .D0(n6209), .S0(n306), .D1(n291), .S1(n308), .D2(
        n298), .S2(n280), .D3(n277), .S3(n310), .Z(n6560) );
  HS65_LS_NAND4ABX3 U15961 ( .A(n4967), .B(n4968), .C(n4969), .D(n4970), .Z(
        n4778) );
  HS65_LS_NAND4ABX3 U15962 ( .A(n4996), .B(n4997), .C(n4998), .D(n4999), .Z(
        n4968) );
  HS65_LS_NOR4ABX2 U15963 ( .A(n4971), .B(n4972), .C(n4973), .D(n4974), .Z(
        n4970) );
  HS65_LS_MX41X4 U15964 ( .D0(n4616), .S0(n483), .D1(n468), .S1(n485), .D2(
        n475), .S2(n457), .D3(n454), .S3(n487), .Z(n4967) );
  HS65_LS_NAND4ABX3 U15965 ( .A(n4913), .B(n4914), .C(n4915), .D(n4916), .Z(
        n4739) );
  HS65_LS_NAND4ABX3 U15966 ( .A(n4942), .B(n4943), .C(n4944), .D(n4945), .Z(
        n4914) );
  HS65_LS_NOR4ABX2 U15967 ( .A(n4917), .B(n4918), .C(n4919), .D(n4920), .Z(
        n4916) );
  HS65_LS_MX41X4 U15968 ( .D0(n4591), .S0(n264), .D1(n249), .S1(n266), .D2(
        n256), .S2(n238), .D3(n235), .S3(n268), .Z(n4913) );
  HS65_LS_NAND4ABX3 U15969 ( .A(n4837), .B(n4838), .C(n4839), .D(n4840), .Z(
        n4631) );
  HS65_LS_NAND4ABX3 U15970 ( .A(n4868), .B(n4869), .C(n4870), .D(n4871), .Z(
        n4838) );
  HS65_LS_NOR4ABX2 U15971 ( .A(n4841), .B(n4842), .C(n4843), .D(n4844), .Z(
        n4840) );
  HS65_LS_MX41X4 U15972 ( .D0(n4531), .S0(n701), .D1(n676), .S1(n707), .D2(
        n709), .S2(n684), .D3(n688), .S3(n704), .Z(n4837) );
  HS65_LS_NAND4ABX3 U15973 ( .A(n6430), .B(n6431), .C(n6432), .D(n6433), .Z(
        n6224) );
  HS65_LS_NAND4ABX3 U15974 ( .A(n6461), .B(n6462), .C(n6463), .D(n6464), .Z(
        n6431) );
  HS65_LS_NOR4ABX2 U15975 ( .A(n6434), .B(n6435), .C(n6436), .D(n6437), .Z(
        n6433) );
  HS65_LS_MX41X4 U15976 ( .D0(n6124), .S0(n519), .D1(n494), .S1(n525), .D2(
        n527), .S2(n502), .D3(n506), .S3(n522), .Z(n6430) );
  HS65_LS_NAND4ABX3 U15977 ( .A(n4697), .B(n4698), .C(n4699), .D(n4700), .Z(
        n4554) );
  HS65_LS_NAND4ABX3 U15978 ( .A(n4728), .B(n4729), .C(n4730), .D(n4731), .Z(
        n4698) );
  HS65_LS_MX41X4 U15979 ( .D0(n4491), .S0(n37), .D1(n11), .S1(n43), .D2(n45), 
        .S2(n20), .D3(n40), .S3(n24), .Z(n4697) );
  HS65_LS_NOR4ABX2 U15980 ( .A(n4701), .B(n4702), .C(n4703), .D(n4704), .Z(
        n4700) );
  HS65_LS_NAND4ABX3 U15981 ( .A(n6290), .B(n6291), .C(n6292), .D(n6293), .Z(
        n6147) );
  HS65_LS_NAND4ABX3 U15982 ( .A(n6321), .B(n6322), .C(n6323), .D(n6324), .Z(
        n6291) );
  HS65_LS_MX41X4 U15983 ( .D0(n6084), .S0(n563), .D1(n537), .S1(n569), .D2(
        n571), .S2(n546), .D3(n566), .S3(n550), .Z(n6290) );
  HS65_LS_NOR4ABX2 U15984 ( .A(n6294), .B(n6295), .C(n6296), .D(n6297), .Z(
        n6293) );
  HS65_LS_NOR4ABX2 U15985 ( .A(n3949), .B(n3950), .C(n3951), .D(n3952), .Z(
        n3948) );
  HS65_LS_OAI212X3 U15986 ( .A(n3353), .B(n3778), .C(n3148), .D(n2895), .E(
        n2889), .Z(n3951) );
  HS65_LS_IVX2 U15987 ( .A(n7932), .Z(n127) );
  HS65_LS_IVX2 U15988 ( .A(n7833), .Z(n614) );
  HS65_LS_NOR2X2 U15989 ( .A(n7639), .B(n8699), .Z(n8416) );
  HS65_LS_NOR2X2 U15990 ( .A(n7667), .B(n8787), .Z(n8476) );
  HS65_LS_IVX2 U15991 ( .A(n3282), .Z(n149) );
  HS65_LS_NOR4ABX2 U15992 ( .A(n3885), .B(n3886), .C(n3887), .D(n3888), .Z(
        n3367) );
  HS65_LS_NOR3X1 U15993 ( .A(n3897), .B(n3898), .C(n3899), .Z(n3886) );
  HS65_LS_NAND4ABX3 U15994 ( .A(n3889), .B(n2858), .C(n3890), .D(n3891), .Z(
        n3888) );
  HS65_LS_OAI212X3 U15995 ( .A(n3892), .B(n3893), .C(n3894), .D(n3895), .E(
        n3896), .Z(n3887) );
  HS65_LS_IVX2 U15996 ( .A(n1129), .Z(n855) );
  HS65_LS_IVX2 U15997 ( .A(n1881), .Z(n773) );
  HS65_LS_IVX2 U15998 ( .A(n1505), .Z(n814) );
  HS65_LS_IVX2 U15999 ( .A(n2257), .Z(n896) );
  HS65_LS_NOR2X2 U16000 ( .A(n7964), .B(n8051), .Z(n8536) );
  HS65_LS_IVX2 U16001 ( .A(n7861), .Z(n377) );
  HS65_LS_IVX2 U16002 ( .A(n7963), .Z(n326) );
  HS65_LS_NOR2X2 U16003 ( .A(n3776), .B(n3778), .Z(n3697) );
  HS65_LS_NOR2X2 U16004 ( .A(n8412), .B(n7645), .Z(n8166) );
  HS65_LS_NOR2X2 U16005 ( .A(n8472), .B(n7673), .Z(n8198) );
  HS65_LS_NOR4ABX2 U16006 ( .A(n8371), .B(n8372), .C(n8373), .D(n8374), .Z(
        n7948) );
  HS65_LS_OAI212X3 U16007 ( .A(n8378), .B(n8379), .C(n8040), .D(n8335), .E(
        n8380), .Z(n8373) );
  HS65_LS_NAND3X2 U16008 ( .A(n8375), .B(n8376), .C(n8377), .Z(n8374) );
  HS65_LS_AOI222X2 U16009 ( .A(n335), .B(n353), .C(n357), .D(n334), .E(n337), 
        .F(n348), .Z(n8371) );
  HS65_LS_NOR4ABX2 U16010 ( .A(n8497), .B(n8498), .C(n7766), .D(n8499), .Z(
        n8496) );
  HS65_LS_OA212X4 U16011 ( .A(n7761), .B(n8130), .C(n7872), .D(n8019), .E(
        n8505), .Z(n8498) );
  HS65_LS_NOR4ABX2 U16012 ( .A(n8859), .B(n8860), .C(n7783), .D(n8632), .Z(
        n8858) );
  HS65_LS_OA212X4 U16013 ( .A(n7778), .B(n8326), .C(n7955), .D(n8061), .E(
        n8879), .Z(n8860) );
  HS65_LS_NOR2X2 U16014 ( .A(n3536), .B(n3486), .Z(n3456) );
  HS65_LS_NOR2X2 U16015 ( .A(n6339), .B(n6050), .Z(n6900) );
  HS65_LS_NOR2X2 U16016 ( .A(n6232), .B(n6428), .Z(n6784) );
  HS65_LS_NOR2X2 U16017 ( .A(n4639), .B(n4835), .Z(n5192) );
  HS65_LS_NOR2X2 U16018 ( .A(n4785), .B(n4503), .Z(n5423) );
  HS65_LS_NOR2X2 U16019 ( .A(n6378), .B(n6096), .Z(n7015) );
  HS65_LS_NOR2X2 U16020 ( .A(n4746), .B(n4457), .Z(n5308) );
  HS65_LS_IVX2 U16021 ( .A(n7954), .Z(n346) );
  HS65_LS_NAND2X2 U16022 ( .A(n2314), .B(n2263), .Z(n2493) );
  HS65_LS_NAND2X2 U16023 ( .A(n1562), .B(n1511), .Z(n1741) );
  HS65_LS_NOR2X2 U16024 ( .A(n7857), .B(n8019), .Z(n8021) );
  HS65_LS_NOR2X2 U16025 ( .A(n8136), .B(n8019), .Z(n8028) );
  HS65_LS_NOR2X2 U16026 ( .A(n7959), .B(n8061), .Z(n8063) );
  HS65_LS_NAND3X2 U16027 ( .A(n6262), .B(n7116), .C(n6168), .Z(n7119) );
  HS65_LS_NAND3X2 U16028 ( .A(n4669), .B(n5524), .C(n4575), .Z(n5527) );
  HS65_LS_CBI4I1X3 U16029 ( .A(n1154), .B(n1155), .C(n1156), .D(n1157), .Z(
        n1144) );
  HS65_LS_OAI21X2 U16030 ( .A(n854), .B(n869), .C(n882), .Z(n1157) );
  HS65_LS_CBI4I1X3 U16031 ( .A(n1906), .B(n1907), .C(n1908), .D(n1909), .Z(
        n1896) );
  HS65_LS_OAI21X2 U16032 ( .A(n772), .B(n787), .C(n800), .Z(n1909) );
  HS65_LS_NOR2X2 U16033 ( .A(n6872), .B(n7191), .Z(n6923) );
  HS65_LS_NOR2X2 U16034 ( .A(n5280), .B(n5599), .Z(n5331) );
  HS65_LS_NOR2X2 U16035 ( .A(n5395), .B(n5626), .Z(n5446) );
  HS65_LS_NOR2X2 U16036 ( .A(n6987), .B(n7218), .Z(n7038) );
  HS65_LS_NOR2X2 U16037 ( .A(n6755), .B(n7174), .Z(n6807) );
  HS65_LS_NOR2X2 U16038 ( .A(n5163), .B(n5582), .Z(n5215) );
  HS65_LS_IVX2 U16039 ( .A(n3329), .Z(n640) );
  HS65_LS_NOR2X2 U16040 ( .A(n1376), .B(n1312), .Z(n1362) );
  HS65_LS_NOR2X2 U16041 ( .A(n2504), .B(n2440), .Z(n2490) );
  HS65_LS_NOR2X2 U16042 ( .A(n2128), .B(n2064), .Z(n2114) );
  HS65_LS_NOR2X2 U16043 ( .A(n1752), .B(n1688), .Z(n1738) );
  HS65_LS_IVX2 U16044 ( .A(n8663), .Z(n402) );
  HS65_LS_CBI4I1X3 U16045 ( .A(n1686), .B(n1503), .C(n1576), .D(n1806), .Z(
        n1784) );
  HS65_LS_AO12X4 U16046 ( .A(n1775), .B(n1535), .C(n1562), .Z(n1806) );
  HS65_LS_CBI4I1X3 U16047 ( .A(n2438), .B(n2255), .C(n2328), .D(n2558), .Z(
        n2536) );
  HS65_LS_AO12X4 U16048 ( .A(n2527), .B(n2287), .C(n2314), .Z(n2558) );
  HS65_LS_NOR2X2 U16049 ( .A(n3043), .B(n3281), .Z(n3271) );
  HS65_LS_NOR2X2 U16050 ( .A(n3043), .B(n2924), .Z(n3580) );
  HS65_LS_IVX2 U16051 ( .A(n3214), .Z(n431) );
  HS65_LS_IVX2 U16052 ( .A(n4720), .Z(n25) );
  HS65_LS_IVX2 U16053 ( .A(n6313), .Z(n551) );
  HS65_LS_CBI4I1X3 U16054 ( .A(n1310), .B(n1127), .C(n1200), .D(n1430), .Z(
        n1408) );
  HS65_LS_AO12X4 U16055 ( .A(n1399), .B(n1159), .C(n1186), .Z(n1430) );
  HS65_LS_NOR2X2 U16056 ( .A(n2944), .B(n3133), .Z(n3482) );
  HS65_LS_IVX2 U16057 ( .A(n4859), .Z(n689) );
  HS65_LS_IVX2 U16058 ( .A(n4989), .Z(n455) );
  HS65_LS_IVX2 U16059 ( .A(n6582), .Z(n278) );
  HS65_LS_IVX2 U16060 ( .A(n6528), .Z(n57) );
  HS65_LS_IVX2 U16061 ( .A(n6452), .Z(n507) );
  HS65_LS_IVX2 U16062 ( .A(n4935), .Z(n236) );
  HS65_LS_NAND2X2 U16063 ( .A(n1186), .B(n1135), .Z(n1365) );
  HS65_LS_NAND2X2 U16064 ( .A(n1938), .B(n1887), .Z(n2117) );
  HS65_LS_CBI4I1X3 U16065 ( .A(n2062), .B(n1879), .C(n1952), .D(n2182), .Z(
        n2160) );
  HS65_LS_AO12X4 U16066 ( .A(n2151), .B(n1911), .C(n1938), .Z(n2182) );
  HS65_LS_NOR2X2 U16067 ( .A(n3391), .B(n3214), .Z(n3191) );
  HS65_LS_NOR3AX2 U16068 ( .A(n8631), .B(n8895), .C(n8867), .Z(n8889) );
  HS65_LS_OAI21X2 U16069 ( .A(n8045), .B(n8061), .C(n8879), .Z(n8895) );
  HS65_LS_IVX2 U16070 ( .A(n3065), .Z(n182) );
  HS65_LS_IVX2 U16071 ( .A(n3174), .Z(n663) );
  HS65_LS_IVX2 U16072 ( .A(n7645), .Z(n625) );
  HS65_LS_IVX2 U16073 ( .A(n7673), .Z(n138) );
  HS65_LS_NAND2X2 U16074 ( .A(n7777), .B(n7963), .Z(n7775) );
  HS65_LS_NAND2X2 U16075 ( .A(n7760), .B(n7861), .Z(n7758) );
  HS65_LS_IVX2 U16076 ( .A(n3007), .Z(n413) );
  HS65_LS_NOR4ABX2 U16077 ( .A(n3527), .B(n3528), .C(n3529), .D(n3530), .Z(
        n3076) );
  HS65_LS_NOR3X1 U16078 ( .A(n3540), .B(n3541), .C(n3542), .Z(n3528) );
  HS65_LS_OAI212X3 U16079 ( .A(n3535), .B(n3536), .C(n3537), .D(n3538), .E(
        n3539), .Z(n3529) );
  HS65_LS_NAND4ABX3 U16080 ( .A(n3531), .B(n3532), .C(n3533), .D(n3534), .Z(
        n3530) );
  HS65_LS_NOR4ABX2 U16081 ( .A(n3768), .B(n3769), .C(n3770), .D(n3771), .Z(
        n3305) );
  HS65_LS_NOR3X1 U16082 ( .A(n3780), .B(n3781), .C(n3782), .Z(n3769) );
  HS65_LS_OAI212X3 U16083 ( .A(n3775), .B(n3776), .C(n3777), .D(n3778), .E(
        n3779), .Z(n3770) );
  HS65_LS_NAND4ABX3 U16084 ( .A(n3772), .B(n2903), .C(n3773), .D(n3774), .Z(
        n3771) );
  HS65_LS_NOR4ABX2 U16085 ( .A(n8306), .B(n8307), .C(n8308), .D(n8309), .Z(
        n8082) );
  HS65_LS_NOR3X1 U16086 ( .A(n8318), .B(n8319), .C(n8320), .Z(n8307) );
  HS65_LS_NAND4ABX3 U16087 ( .A(n8310), .B(n8311), .C(n8312), .D(n8313), .Z(
        n8309) );
  HS65_LS_OAI212X3 U16088 ( .A(n8314), .B(n8315), .C(n8316), .D(n7761), .E(
        n8317), .Z(n8308) );
  HS65_LS_NAND4ABX3 U16089 ( .A(n1231), .B(n1232), .C(n1233), .D(n1234), .Z(
        n1151) );
  HS65_LS_OAI222X2 U16090 ( .A(n1129), .B(n1155), .C(n1173), .D(n1243), .E(
        n1121), .F(n1127), .Z(n1232) );
  HS65_LS_NOR4ABX2 U16091 ( .A(n1235), .B(n1236), .C(n1237), .D(n1238), .Z(
        n1234) );
  HS65_LS_NOR4ABX2 U16092 ( .A(n1239), .B(n1240), .C(n1241), .D(n1242), .Z(
        n1233) );
  HS65_LS_NAND4ABX3 U16093 ( .A(n2359), .B(n2360), .C(n2361), .D(n2362), .Z(
        n2279) );
  HS65_LS_OAI222X2 U16094 ( .A(n2257), .B(n2283), .C(n2301), .D(n2371), .E(
        n2249), .F(n2255), .Z(n2360) );
  HS65_LS_NOR4ABX2 U16095 ( .A(n2363), .B(n2364), .C(n2365), .D(n2366), .Z(
        n2362) );
  HS65_LS_NAND3AX3 U16096 ( .A(n2372), .B(n2373), .C(n2374), .Z(n2359) );
  HS65_LS_NAND4ABX3 U16097 ( .A(n1983), .B(n1984), .C(n1985), .D(n1986), .Z(
        n1903) );
  HS65_LS_OAI222X2 U16098 ( .A(n1881), .B(n1907), .C(n1925), .D(n1995), .E(
        n1873), .F(n1879), .Z(n1984) );
  HS65_LS_NOR4ABX2 U16099 ( .A(n1987), .B(n1988), .C(n1989), .D(n1990), .Z(
        n1986) );
  HS65_LS_NOR4ABX2 U16100 ( .A(n1991), .B(n1992), .C(n1993), .D(n1994), .Z(
        n1985) );
  HS65_LS_NAND4ABX3 U16101 ( .A(n1607), .B(n1608), .C(n1609), .D(n1610), .Z(
        n1527) );
  HS65_LS_OAI222X2 U16102 ( .A(n1505), .B(n1531), .C(n1549), .D(n1619), .E(
        n1497), .F(n1503), .Z(n1608) );
  HS65_LS_NOR4ABX2 U16103 ( .A(n1611), .B(n1612), .C(n1613), .D(n1614), .Z(
        n1610) );
  HS65_LS_NAND3AX3 U16104 ( .A(n1620), .B(n1621), .C(n1622), .Z(n1607) );
  HS65_LS_NOR2X2 U16105 ( .A(n2985), .B(n2887), .Z(n3343) );
  HS65_LS_NOR2X2 U16106 ( .A(n3146), .B(n3359), .Z(n3723) );
  HS65_LS_IVX2 U16107 ( .A(n3173), .Z(n655) );
  HS65_LS_NAND4ABX3 U16108 ( .A(n4134), .B(n4135), .C(n4136), .D(n4137), .Z(
        n3927) );
  HS65_LS_NOR4ABX2 U16109 ( .A(n3638), .B(n3663), .C(n3620), .D(n3265), .Z(
        n4136) );
  HS65_LS_CBI4I1X3 U16110 ( .A(n3067), .B(n3297), .C(n2925), .D(n3561), .Z(
        n4134) );
  HS65_LS_CBI4I1X3 U16111 ( .A(n173), .B(n3066), .C(n3063), .D(n4166), .Z(
        n4135) );
  HS65_LS_NAND2X2 U16112 ( .A(n8220), .B(n7862), .Z(n8218) );
  HS65_LS_NAND4ABX3 U16113 ( .A(n2143), .B(n2144), .C(n2145), .D(n2146), .Z(
        n1876) );
  HS65_LS_CBI4I1X3 U16114 ( .A(n1873), .B(n1966), .C(n1908), .D(n1988), .Z(
        n2143) );
  HS65_LS_NOR4ABX2 U16115 ( .A(n2032), .B(n2054), .C(n2075), .D(n2098), .Z(
        n2145) );
  HS65_LS_CBI4I1X3 U16116 ( .A(n779), .B(n2153), .C(n1886), .D(n2154), .Z(
        n2144) );
  HS65_LS_NAND4ABX3 U16117 ( .A(n1391), .B(n1392), .C(n1393), .D(n1394), .Z(
        n1124) );
  HS65_LS_CBI4I1X3 U16118 ( .A(n1121), .B(n1214), .C(n1156), .D(n1236), .Z(
        n1391) );
  HS65_LS_NOR4ABX2 U16119 ( .A(n1280), .B(n1302), .C(n1323), .D(n1346), .Z(
        n1393) );
  HS65_LS_CBI4I1X3 U16120 ( .A(n861), .B(n1401), .C(n1134), .D(n1402), .Z(
        n1392) );
  HS65_LS_NAND4ABX3 U16121 ( .A(n1767), .B(n1768), .C(n1769), .D(n1770), .Z(
        n1500) );
  HS65_LS_CBI4I1X3 U16122 ( .A(n1497), .B(n1590), .C(n1532), .D(n1612), .Z(
        n1767) );
  HS65_LS_NOR4ABX2 U16123 ( .A(n1656), .B(n1678), .C(n1699), .D(n1722), .Z(
        n1769) );
  HS65_LS_CBI4I1X3 U16124 ( .A(n820), .B(n1777), .C(n1510), .D(n1778), .Z(
        n1768) );
  HS65_LS_NAND4ABX3 U16125 ( .A(n2519), .B(n2520), .C(n2521), .D(n2522), .Z(
        n2252) );
  HS65_LS_CBI4I1X3 U16126 ( .A(n2249), .B(n2342), .C(n2284), .D(n2364), .Z(
        n2519) );
  HS65_LS_NOR4ABX2 U16127 ( .A(n2408), .B(n2430), .C(n2451), .D(n2474), .Z(
        n2521) );
  HS65_LS_CBI4I1X3 U16128 ( .A(n902), .B(n2529), .C(n2262), .D(n2530), .Z(
        n2520) );
  HS65_LS_NOR2X2 U16129 ( .A(n7663), .B(n8787), .Z(n8826) );
  HS65_LS_NOR2X2 U16130 ( .A(n7635), .B(n8699), .Z(n8738) );
  HS65_LS_IVX2 U16131 ( .A(n8639), .Z(n343) );
  HS65_LS_IVX2 U16132 ( .A(n1243), .Z(n884) );
  HS65_LS_IVX2 U16133 ( .A(n1995), .Z(n802) );
  HS65_LS_IVX2 U16134 ( .A(n2371), .Z(n925) );
  HS65_LS_IVX2 U16135 ( .A(n1619), .Z(n843) );
  HS65_LS_NOR2X2 U16136 ( .A(n2893), .B(n3174), .Z(n3782) );
  HS65_LS_IVX2 U16137 ( .A(n8018), .Z(n398) );
  HS65_LS_IVX2 U16138 ( .A(n8060), .Z(n351) );
  HS65_LS_NOR2X2 U16139 ( .A(n3329), .B(n3173), .Z(n3150) );
  HS65_LS_NAND2X2 U16140 ( .A(n7670), .B(n7885), .Z(n7733) );
  HS65_LS_NAND2X2 U16141 ( .A(n7642), .B(n7846), .Z(n7695) );
  HS65_LS_NAND2X2 U16142 ( .A(n3538), .B(n3905), .Z(n3451) );
  HS65_LS_NAND2X2 U16143 ( .A(n3778), .B(n2900), .Z(n3695) );
  HS65_LS_IVX2 U16144 ( .A(n7735), .Z(n111) );
  HS65_LS_IVX2 U16145 ( .A(n7697), .Z(n598) );
  HS65_LS_IVX2 U16146 ( .A(n8136), .Z(n380) );
  HS65_LS_NAND2X2 U16147 ( .A(n7761), .B(n7870), .Z(n8217) );
  HS65_LS_IVX2 U16148 ( .A(n2842), .Z(n445) );
  HS65_LS_IVX2 U16149 ( .A(n7858), .Z(n381) );
  HS65_LS_IVX2 U16150 ( .A(n7960), .Z(n332) );
  HS65_LS_IVX2 U16151 ( .A(n1155), .Z(n880) );
  HS65_LS_IVX2 U16152 ( .A(n1907), .Z(n798) );
  HS65_LS_AOI12X2 U16153 ( .A(n2960), .B(n3538), .C(n2961), .Z(n4183) );
  HS65_LS_IVX2 U16154 ( .A(n2283), .Z(n921) );
  HS65_LS_IVX2 U16155 ( .A(n1531), .Z(n839) );
  HS65_LS_NAND2X2 U16156 ( .A(n46), .B(n4491), .Z(n4711) );
  HS65_LS_NAND2X2 U16157 ( .A(n572), .B(n6084), .Z(n6304) );
  HS65_LS_NOR2X2 U16158 ( .A(n8046), .B(n8379), .Z(n8598) );
  HS65_LS_IVX2 U16159 ( .A(n8069), .Z(n330) );
  HS65_LS_NOR2X2 U16160 ( .A(n2371), .B(n2527), .Z(n2303) );
  HS65_LS_NOR2X2 U16161 ( .A(n1619), .B(n1775), .Z(n1551) );
  HS65_LS_IVX2 U16162 ( .A(n3359), .Z(n637) );
  HS65_LS_IVX2 U16163 ( .A(n3421), .Z(n414) );
  HS65_LS_NAND2X2 U16164 ( .A(n8220), .B(n8030), .Z(n8250) );
  HS65_LS_NOR2X2 U16165 ( .A(n7959), .B(n8379), .Z(n8382) );
  HS65_LS_NOR2X2 U16166 ( .A(n4559), .B(n4676), .Z(n5035) );
  HS65_LS_NOR2X2 U16167 ( .A(n6152), .B(n6269), .Z(n6628) );
  HS65_LS_NAND2X2 U16168 ( .A(n3454), .B(n2878), .Z(n3452) );
  HS65_LS_NAND2X2 U16169 ( .A(n76), .B(n6184), .Z(n6520) );
  HS65_LS_NAND2X2 U16170 ( .A(n297), .B(n6209), .Z(n6574) );
  HS65_LS_NAND2X2 U16171 ( .A(n474), .B(n4616), .Z(n4981) );
  HS65_LS_NAND2X2 U16172 ( .A(n255), .B(n4591), .Z(n4927) );
  HS65_LS_NAND2X2 U16173 ( .A(n710), .B(n4531), .Z(n4851) );
  HS65_LS_NAND2X2 U16174 ( .A(n528), .B(n6124), .Z(n6444) );
  HS65_LS_NOR2X2 U16175 ( .A(n1243), .B(n1399), .Z(n1175) );
  HS65_LS_NOR2X2 U16176 ( .A(n4783), .B(n5008), .Z(n5390) );
  HS65_LS_NOR2X2 U16177 ( .A(n4744), .B(n4894), .Z(n5275) );
  HS65_LS_NOR2X2 U16178 ( .A(n4637), .B(n4880), .Z(n5158) );
  HS65_LS_NOR2X2 U16179 ( .A(n6376), .B(n6601), .Z(n6982) );
  HS65_LS_NOR2X2 U16180 ( .A(n6230), .B(n6473), .Z(n6750) );
  HS65_LS_NOR2X2 U16181 ( .A(n6337), .B(n6487), .Z(n6867) );
  HS65_LS_IVX2 U16182 ( .A(n4722), .Z(n40) );
  HS65_LS_IVX2 U16183 ( .A(n6315), .Z(n566) );
  HS65_LS_IVX2 U16184 ( .A(n2971), .Z(n228) );
  HS65_LS_NAND2X2 U16185 ( .A(n7931), .B(n7880), .Z(n8824) );
  HS65_LS_NAND2X2 U16186 ( .A(n7832), .B(n7817), .Z(n8736) );
  HS65_LS_NAND2X2 U16187 ( .A(n608), .B(n7709), .Z(n8407) );
  HS65_LS_NAND2X2 U16188 ( .A(n121), .B(n7747), .Z(n8467) );
  HS65_LS_IVX2 U16189 ( .A(n7779), .Z(n357) );
  HS65_LS_IVX2 U16190 ( .A(n8051), .Z(n352) );
  HS65_LS_NOR2X2 U16191 ( .A(n1995), .B(n2151), .Z(n1927) );
  HS65_LS_NOR2X2 U16192 ( .A(n6288), .B(n6634), .Z(n6656) );
  HS65_LS_NOR2X2 U16193 ( .A(n4695), .B(n5041), .Z(n5063) );
  HS65_LS_IVX2 U16194 ( .A(n2854), .Z(n424) );
  HS65_LS_IVX2 U16195 ( .A(n7762), .Z(n393) );
  HS65_LS_NAND3X2 U16196 ( .A(n3065), .B(n3290), .C(n3051), .Z(n4004) );
  HS65_LS_NOR3AX2 U16197 ( .A(n8650), .B(n8955), .C(n8658), .Z(n8949) );
  HS65_LS_OAI21X2 U16198 ( .A(n8003), .B(n8019), .C(n8505), .Z(n8955) );
  HS65_LS_NAND2X2 U16199 ( .A(n3599), .B(n2928), .Z(n3597) );
  HS65_LS_NAND2X2 U16200 ( .A(n555), .B(n6084), .Z(n6625) );
  HS65_LS_NAND2X2 U16201 ( .A(n29), .B(n4491), .Z(n5032) );
  HS65_LS_IVX2 U16202 ( .A(n8186), .Z(n110) );
  HS65_LS_IVX2 U16203 ( .A(n8154), .Z(n597) );
  HS65_LS_IVX2 U16204 ( .A(n3004), .Z(n417) );
  HS65_LS_NOR2X2 U16205 ( .A(n8019), .B(n7861), .Z(n8245) );
  HS65_LS_NOR2X2 U16206 ( .A(n8061), .B(n7963), .Z(n8549) );
  HS65_LS_NOR2X2 U16207 ( .A(n7960), .B(n8639), .Z(n8048) );
  HS65_LS_NOR2X2 U16208 ( .A(n3585), .B(n3281), .Z(n3592) );
  HS65_LS_NOR2X2 U16209 ( .A(n7963), .B(n8639), .Z(n8329) );
  HS65_LS_OAI21X2 U16210 ( .A(n6065), .B(n6051), .C(n6491), .Z(n6490) );
  HS65_LS_OAI21X2 U16211 ( .A(n6111), .B(n6097), .C(n6545), .Z(n6544) );
  HS65_LS_OAI21X2 U16212 ( .A(n4472), .B(n4458), .C(n4898), .Z(n4897) );
  HS65_LS_OAI21X2 U16213 ( .A(n4518), .B(n4504), .C(n4952), .Z(n4951) );
  HS65_LS_OAI21X2 U16214 ( .A(n4533), .B(n4820), .C(n4821), .Z(n4819) );
  HS65_LS_OAI21X2 U16215 ( .A(n6126), .B(n6413), .C(n6414), .Z(n6412) );
  HS65_LS_IVX2 U16216 ( .A(n7886), .Z(n132) );
  HS65_LS_IVX2 U16217 ( .A(n7847), .Z(n619) );
  HS65_LS_IVX2 U16218 ( .A(n7634), .Z(n591) );
  HS65_LS_IVX2 U16219 ( .A(n7662), .Z(n104) );
  HS65_LS_NAND2X2 U16220 ( .A(n81), .B(n6184), .Z(n6862) );
  HS65_LS_NAND2X2 U16221 ( .A(n260), .B(n4591), .Z(n5270) );
  HS65_LS_NAND2X2 U16222 ( .A(n479), .B(n4616), .Z(n5385) );
  HS65_LS_NAND2X2 U16223 ( .A(n302), .B(n6209), .Z(n6977) );
  HS65_LS_NAND2X2 U16224 ( .A(n693), .B(n4531), .Z(n5153) );
  HS65_LS_NAND2X2 U16225 ( .A(n511), .B(n6124), .Z(n6745) );
  HS65_LS_IVX2 U16226 ( .A(n3263), .Z(n156) );
  HS65_LS_NAND3X2 U16227 ( .A(n6481), .B(n7136), .C(n6352), .Z(n7211) );
  HS65_LS_NAND3X2 U16228 ( .A(n5002), .B(n5565), .C(n4798), .Z(n5646) );
  HS65_LS_NAND3X2 U16229 ( .A(n6595), .B(n7157), .C(n6391), .Z(n7238) );
  HS65_LS_NAND3X2 U16230 ( .A(n4888), .B(n5544), .C(n4759), .Z(n5619) );
  HS65_LS_NAND3X2 U16231 ( .A(n4874), .B(n5589), .C(n4652), .Z(n5592) );
  HS65_LS_NAND3X2 U16232 ( .A(n6467), .B(n7181), .C(n6245), .Z(n7184) );
  HS65_LS_IVX2 U16233 ( .A(n2924), .Z(n155) );
  HS65_LS_NOR2X2 U16234 ( .A(n3127), .B(n3133), .Z(n3532) );
  HS65_LS_IVX2 U16235 ( .A(n6314), .Z(n552) );
  HS65_LS_IVX2 U16236 ( .A(n4721), .Z(n26) );
  HS65_LS_IVX2 U16237 ( .A(n4861), .Z(n690) );
  HS65_LS_IVX2 U16238 ( .A(n4990), .Z(n456) );
  HS65_LS_IVX2 U16239 ( .A(n6583), .Z(n279) );
  HS65_LS_IVX2 U16240 ( .A(n6529), .Z(n58) );
  HS65_LS_IVX2 U16241 ( .A(n6454), .Z(n508) );
  HS65_LS_IVX2 U16242 ( .A(n4936), .Z(n237) );
  HS65_LS_NOR2X2 U16243 ( .A(n3415), .B(n3421), .Z(n2858) );
  HS65_LS_NOR2X2 U16244 ( .A(n8192), .B(n7673), .Z(n8833) );
  HS65_LS_NOR2X2 U16245 ( .A(n8160), .B(n7645), .Z(n8745) );
  HS65_LS_NAND2X2 U16246 ( .A(n7832), .B(n8159), .Z(n8688) );
  HS65_LS_NAND2X2 U16247 ( .A(n7931), .B(n8191), .Z(n8776) );
  HS65_LS_NOR2X2 U16248 ( .A(n8119), .B(n7760), .Z(n8022) );
  HS65_LS_NOR2X2 U16249 ( .A(n6634), .B(n6154), .Z(n6166) );
  HS65_LS_NOR2X2 U16250 ( .A(n5041), .B(n4561), .Z(n4573) );
  HS65_LS_OAI21X2 U16251 ( .A(n3064), .B(n3067), .C(n4090), .Z(n4116) );
  HS65_LS_NAND2X2 U16252 ( .A(n623), .B(n7709), .Z(n8696) );
  HS65_LS_NAND2X2 U16253 ( .A(n136), .B(n7747), .Z(n8784) );
  HS65_LS_NOR2X2 U16254 ( .A(n2848), .B(n3214), .Z(n3791) );
  HS65_LS_IVX2 U16255 ( .A(n1498), .Z(n824) );
  HS65_LS_IVX2 U16256 ( .A(n2250), .Z(n906) );
  HS65_LS_IVX2 U16257 ( .A(n3391), .Z(n416) );
  HS65_LS_OAI21X2 U16258 ( .A(n7847), .B(n7686), .C(n8390), .Z(n8389) );
  HS65_LS_OAI21X2 U16259 ( .A(n7886), .B(n7724), .C(n8450), .Z(n8449) );
  HS65_LS_OAI21X2 U16260 ( .A(n7893), .B(n7724), .C(n7737), .Z(n7892) );
  HS65_LS_OAI21X2 U16261 ( .A(n7793), .B(n7686), .C(n7699), .Z(n7792) );
  HS65_LS_NAND2X2 U16262 ( .A(n3599), .B(n3263), .Z(n3609) );
  HS65_LS_OAI21X2 U16263 ( .A(n3236), .B(n3067), .C(n3237), .Z(n3235) );
  HS65_LS_NAND2X2 U16264 ( .A(n2281), .B(n2256), .Z(n2494) );
  HS65_LS_NAND2X2 U16265 ( .A(n1529), .B(n1504), .Z(n1742) );
  HS65_LS_IVX2 U16266 ( .A(n8030), .Z(n379) );
  HS65_LS_IVX2 U16267 ( .A(n1122), .Z(n865) );
  HS65_LS_IVX2 U16268 ( .A(n1874), .Z(n783) );
  HS65_LS_IVX2 U16269 ( .A(n2874), .Z(n200) );
  HS65_LS_IVX2 U16270 ( .A(n6194), .Z(n62) );
  HS65_LS_IVX2 U16271 ( .A(n4601), .Z(n241) );
  HS65_LS_IVX2 U16272 ( .A(n4613), .Z(n460) );
  HS65_LS_IVX2 U16273 ( .A(n6206), .Z(n283) );
  HS65_LS_IVX2 U16274 ( .A(n6136), .Z(n504) );
  HS65_LS_IVX2 U16275 ( .A(n4543), .Z(n686) );
  HS65_LS_OAI21X2 U16276 ( .A(n3893), .B(n3414), .C(n4300), .Z(n4299) );
  HS65_LS_OAI21X2 U16277 ( .A(n425), .B(n419), .C(n443), .Z(n4300) );
  HS65_LS_IVX2 U16278 ( .A(n8159), .Z(n596) );
  HS65_LS_IVX2 U16279 ( .A(n8191), .Z(n109) );
  HS65_LS_NOR2AX3 U16280 ( .A(n6084), .B(n6312), .Z(n6158) );
  HS65_LS_NOR2AX3 U16281 ( .A(n4491), .B(n4719), .Z(n4565) );
  HS65_LS_IVX2 U16282 ( .A(n5008), .Z(n453) );
  HS65_LS_IVX2 U16283 ( .A(n4894), .Z(n234) );
  HS65_LS_IVX2 U16284 ( .A(n6601), .Z(n276) );
  HS65_LS_IVX2 U16285 ( .A(n6487), .Z(n55) );
  HS65_LS_IVX2 U16286 ( .A(n4880), .Z(n687) );
  HS65_LS_IVX2 U16287 ( .A(n6473), .Z(n505) );
  HS65_LS_NOR2X2 U16288 ( .A(n7761), .B(n8018), .Z(n8126) );
  HS65_LS_NOR2AX3 U16289 ( .A(n6184), .B(n6059), .Z(n6342) );
  HS65_LS_NOR2AX3 U16290 ( .A(n4616), .B(n4512), .Z(n4788) );
  HS65_LS_NOR2AX3 U16291 ( .A(n6209), .B(n6105), .Z(n6381) );
  HS65_LS_NOR2AX3 U16292 ( .A(n4591), .B(n4466), .Z(n4749) );
  HS65_LS_NOR2AX3 U16293 ( .A(n4531), .B(n4860), .Z(n4642) );
  HS65_LS_NOR2X2 U16294 ( .A(n7778), .B(n8060), .Z(n8368) );
  HS65_LS_NOR2AX3 U16295 ( .A(n6124), .B(n6453), .Z(n6235) );
  HS65_LS_NAND2X2 U16296 ( .A(n1153), .B(n1128), .Z(n1366) );
  HS65_LS_NAND2X2 U16297 ( .A(n1905), .B(n1880), .Z(n2118) );
  HS65_LS_OAI21X2 U16298 ( .A(n4503), .B(n4504), .C(n4505), .Z(n4502) );
  HS65_LS_OAI21X2 U16299 ( .A(n4457), .B(n4458), .C(n4459), .Z(n4456) );
  HS65_LS_OAI21X2 U16300 ( .A(n6096), .B(n6097), .C(n6098), .Z(n6095) );
  HS65_LS_OAI21X2 U16301 ( .A(n4835), .B(n4820), .C(n5697), .Z(n5771) );
  HS65_LS_OAI21X2 U16302 ( .A(n6428), .B(n6413), .C(n7289), .Z(n7363) );
  HS65_LS_OAI21X2 U16303 ( .A(n6050), .B(n6051), .C(n6052), .Z(n6049) );
  HS65_LS_NOR2X2 U16304 ( .A(n6872), .B(n6338), .Z(n6350) );
  HS65_LS_NOR2X2 U16305 ( .A(n5395), .B(n4784), .Z(n4796) );
  HS65_LS_NOR2X2 U16306 ( .A(n6987), .B(n6377), .Z(n6389) );
  HS65_LS_NOR2X2 U16307 ( .A(n5280), .B(n4745), .Z(n4757) );
  HS65_LS_NOR2X2 U16308 ( .A(n5163), .B(n4638), .Z(n4650) );
  HS65_LS_NOR2X2 U16309 ( .A(n6755), .B(n6231), .Z(n6243) );
  HS65_LS_NOR2AX3 U16310 ( .A(n6184), .B(n6050), .Z(n6497) );
  HS65_LS_NOR2AX3 U16311 ( .A(n6209), .B(n6096), .Z(n6551) );
  HS65_LS_NOR2AX3 U16312 ( .A(n4591), .B(n4457), .Z(n4904) );
  HS65_LS_NOR2AX3 U16313 ( .A(n4616), .B(n4503), .Z(n4958) );
  HS65_LS_NOR2AX3 U16314 ( .A(n4531), .B(n4835), .Z(n4827) );
  HS65_LS_NOR2AX3 U16315 ( .A(n6124), .B(n6428), .Z(n6420) );
  HS65_LS_NOR2X2 U16316 ( .A(n2301), .B(n2286), .Z(n2480) );
  HS65_LS_NOR2X2 U16317 ( .A(n1549), .B(n1534), .Z(n1728) );
  HS65_LS_NAND4ABX3 U16318 ( .A(n3250), .B(n3251), .C(n3252), .D(n3253), .Z(
        n2920) );
  HS65_LS_OAI222X2 U16319 ( .A(n3262), .B(n2924), .C(n3044), .D(n3263), .E(
        n3264), .F(n3067), .Z(n3251) );
  HS65_LS_NOR4ABX2 U16320 ( .A(n3254), .B(n3255), .C(n3256), .D(n3257), .Z(
        n3253) );
  HS65_LS_NOR4ABX2 U16321 ( .A(n3258), .B(n3259), .C(n3260), .D(n3261), .Z(
        n3252) );
  HS65_LS_NAND4ABX3 U16322 ( .A(n3088), .B(n3089), .C(n3090), .D(n3091), .Z(
        n2870) );
  HS65_LS_OAI222X2 U16323 ( .A(n3100), .B(n2874), .C(n2946), .D(n3101), .E(
        n2973), .F(n3102), .Z(n3089) );
  HS65_LS_NOR4ABX2 U16324 ( .A(n3096), .B(n3097), .C(n3098), .D(n3099), .Z(
        n3090) );
  HS65_LS_NOR4ABX2 U16325 ( .A(n3092), .B(n3093), .C(n3094), .D(n3095), .Z(
        n3091) );
  HS65_LS_NAND4ABX3 U16326 ( .A(n3379), .B(n3380), .C(n3381), .D(n3382), .Z(
        n3000) );
  HS65_LS_OAI222X2 U16327 ( .A(n2849), .B(n3004), .C(n3189), .D(n3391), .E(
        n2841), .F(n2847), .Z(n3380) );
  HS65_LS_NOR4ABX2 U16328 ( .A(n3383), .B(n3384), .C(n3385), .D(n3386), .Z(
        n3382) );
  HS65_LS_NOR4ABX2 U16329 ( .A(n3387), .B(n3388), .C(n3389), .D(n3390), .Z(
        n3381) );
  HS65_LS_OAI21X2 U16330 ( .A(n4493), .B(n4680), .C(n4681), .Z(n4679) );
  HS65_LS_OAI21X2 U16331 ( .A(n6086), .B(n6273), .C(n6274), .Z(n6272) );
  HS65_LS_NAND4ABX3 U16332 ( .A(n3317), .B(n3318), .C(n3319), .D(n3320), .Z(
        n2982) );
  HS65_LS_OAI222X2 U16333 ( .A(n2894), .B(n2986), .C(n3148), .D(n3329), .E(
        n2886), .F(n2892), .Z(n3318) );
  HS65_LS_NOR4ABX2 U16334 ( .A(n3321), .B(n3322), .C(n3323), .D(n3324), .Z(
        n3320) );
  HS65_LS_NAND3AX3 U16335 ( .A(n3330), .B(n3331), .C(n3332), .Z(n3317) );
  HS65_LS_OAI21X2 U16336 ( .A(n5626), .B(n5001), .C(n5893), .Z(n5892) );
  HS65_LS_OAI21X2 U16337 ( .A(n467), .B(n461), .C(n487), .Z(n5893) );
  HS65_LS_OAI21X2 U16338 ( .A(n5599), .B(n4887), .C(n5834), .Z(n5833) );
  HS65_LS_OAI21X2 U16339 ( .A(n248), .B(n242), .C(n268), .Z(n5834) );
  HS65_LS_OAI21X2 U16340 ( .A(n5582), .B(n4873), .C(n5683), .Z(n5682) );
  HS65_LS_OAI21X2 U16341 ( .A(n677), .B(n679), .C(n704), .Z(n5683) );
  HS65_LS_OAI21X2 U16342 ( .A(n7218), .B(n6594), .C(n7485), .Z(n7484) );
  HS65_LS_OAI21X2 U16343 ( .A(n290), .B(n284), .C(n310), .Z(n7485) );
  HS65_LS_OAI21X2 U16344 ( .A(n7191), .B(n6480), .C(n7426), .Z(n7425) );
  HS65_LS_OAI21X2 U16345 ( .A(n69), .B(n63), .C(n89), .Z(n7426) );
  HS65_LS_OAI21X2 U16346 ( .A(n7174), .B(n6466), .C(n7275), .Z(n7274) );
  HS65_LS_OAI21X2 U16347 ( .A(n495), .B(n497), .C(n522), .Z(n7275) );
  HS65_LS_OAI21X2 U16348 ( .A(n3776), .B(n3352), .C(n4241), .Z(n4240) );
  HS65_LS_OAI21X2 U16349 ( .A(n649), .B(n643), .C(n667), .Z(n4241) );
  HS65_LS_NAND2X2 U16350 ( .A(n3002), .B(n2848), .Z(n3813) );
  HS65_LS_NOR2X2 U16351 ( .A(n1173), .B(n1158), .Z(n1352) );
  HS65_LS_NOR2X2 U16352 ( .A(n1925), .B(n1910), .Z(n2104) );
  HS65_LS_NOR2X2 U16353 ( .A(n3189), .B(n3007), .Z(n3823) );
  HS65_LS_NOR2X2 U16354 ( .A(n8136), .B(n8130), .Z(n8311) );
  HS65_LS_NOR2X2 U16355 ( .A(n7638), .B(n8699), .Z(n8702) );
  HS65_LS_NOR2X2 U16356 ( .A(n7666), .B(n8787), .Z(n8790) );
  HS65_LS_NOR2X2 U16357 ( .A(n2299), .B(n2314), .Z(n2378) );
  HS65_LS_NOR2X2 U16358 ( .A(n1547), .B(n1562), .Z(n1626) );
  HS65_LS_NAND2X2 U16359 ( .A(n2281), .B(n2371), .Z(n2423) );
  HS65_LS_NAND2X2 U16360 ( .A(n1529), .B(n1619), .Z(n1671) );
  HS65_LS_NOR2X2 U16361 ( .A(n2946), .B(n2877), .Z(n3463) );
  HS65_LS_NOR2X2 U16362 ( .A(n3148), .B(n2989), .Z(n3706) );
  HS65_LS_NOR2X2 U16363 ( .A(n8018), .B(n8030), .Z(n8238) );
  HS65_LS_NOR2X2 U16364 ( .A(n3067), .B(n3044), .Z(n3270) );
  HS65_LS_NOR2X2 U16365 ( .A(n8267), .B(n7871), .Z(n8268) );
  HS65_LS_IVX2 U16366 ( .A(n3133), .Z(n198) );
  HS65_LS_NOR2X2 U16367 ( .A(n1171), .B(n1186), .Z(n1250) );
  HS65_LS_NOR2X2 U16368 ( .A(n1923), .B(n1938), .Z(n2002) );
  HS65_LS_NAND4ABX3 U16369 ( .A(n6858), .B(n6859), .C(n6860), .D(n6861), .Z(
        n6330) );
  HS65_LS_NOR4ABX2 U16370 ( .A(n6862), .B(n6863), .C(n6864), .D(n6865), .Z(
        n6861) );
  HS65_LS_OAI212X3 U16371 ( .A(n6869), .B(n6870), .C(n6488), .D(n6057), .E(
        n6871), .Z(n6859) );
  HS65_LS_NOR3AX2 U16372 ( .A(n6866), .B(n6867), .C(n6868), .Z(n6860) );
  HS65_LS_NAND4ABX3 U16373 ( .A(n5266), .B(n5267), .C(n5268), .D(n5269), .Z(
        n4737) );
  HS65_LS_NOR4ABX2 U16374 ( .A(n5270), .B(n5271), .C(n5272), .D(n5273), .Z(
        n5269) );
  HS65_LS_OAI212X3 U16375 ( .A(n5277), .B(n5278), .C(n4895), .D(n4464), .E(
        n5279), .Z(n5267) );
  HS65_LS_NOR3AX2 U16376 ( .A(n5274), .B(n5275), .C(n5276), .Z(n5268) );
  HS65_LS_NAND4ABX3 U16377 ( .A(n5381), .B(n5382), .C(n5383), .D(n5384), .Z(
        n4776) );
  HS65_LS_NOR4ABX2 U16378 ( .A(n5385), .B(n5386), .C(n5387), .D(n5388), .Z(
        n5384) );
  HS65_LS_OAI212X3 U16379 ( .A(n5392), .B(n5393), .C(n5009), .D(n4510), .E(
        n5394), .Z(n5382) );
  HS65_LS_NOR3AX2 U16380 ( .A(n5389), .B(n5390), .C(n5391), .Z(n5383) );
  HS65_LS_NAND4ABX3 U16381 ( .A(n6973), .B(n6974), .C(n6975), .D(n6976), .Z(
        n6369) );
  HS65_LS_NOR4ABX2 U16382 ( .A(n6977), .B(n6978), .C(n6979), .D(n6980), .Z(
        n6976) );
  HS65_LS_OAI212X3 U16383 ( .A(n6984), .B(n6985), .C(n6602), .D(n6103), .E(
        n6986), .Z(n6974) );
  HS65_LS_NOR3AX2 U16384 ( .A(n6981), .B(n6982), .C(n6983), .Z(n6975) );
  HS65_LS_NAND4ABX3 U16385 ( .A(n5149), .B(n5150), .C(n5151), .D(n5152), .Z(
        n4629) );
  HS65_LS_NOR4ABX2 U16386 ( .A(n5153), .B(n5154), .C(n5155), .D(n5156), .Z(
        n5152) );
  HS65_LS_OAI212X3 U16387 ( .A(n5160), .B(n5161), .C(n4881), .D(n4544), .E(
        n5162), .Z(n5150) );
  HS65_LS_NOR3AX2 U16388 ( .A(n5157), .B(n5158), .C(n5159), .Z(n5151) );
  HS65_LS_NAND4ABX3 U16389 ( .A(n6741), .B(n6742), .C(n6743), .D(n6744), .Z(
        n6222) );
  HS65_LS_NOR4ABX2 U16390 ( .A(n6745), .B(n6746), .C(n6747), .D(n6748), .Z(
        n6744) );
  HS65_LS_OAI212X3 U16391 ( .A(n6752), .B(n6753), .C(n6474), .D(n6137), .E(
        n6754), .Z(n6742) );
  HS65_LS_NOR3AX2 U16392 ( .A(n6749), .B(n6750), .C(n6751), .Z(n6743) );
  HS65_LS_NOR2X2 U16393 ( .A(n1504), .B(n1775), .Z(n1650) );
  HS65_LS_NOR2X2 U16394 ( .A(n2256), .B(n2527), .Z(n2402) );
  HS65_LS_NOR2X2 U16395 ( .A(n8332), .B(n8326), .Z(n8538) );
  HS65_LS_NAND2X2 U16396 ( .A(n1153), .B(n1243), .Z(n1295) );
  HS65_LS_NAND2X2 U16397 ( .A(n1905), .B(n1995), .Z(n2047) );
  HS65_LS_NAND4ABX3 U16398 ( .A(n6620), .B(n6621), .C(n6622), .D(n6623), .Z(
        n6145) );
  HS65_LS_NOR3X1 U16399 ( .A(n6628), .B(n6629), .C(n6630), .Z(n6622) );
  HS65_LS_NOR4ABX2 U16400 ( .A(n6624), .B(n6625), .C(n6626), .D(n6627), .Z(
        n6623) );
  HS65_LS_OAI212X3 U16401 ( .A(n6631), .B(n6632), .C(n6270), .D(n6081), .E(
        n6633), .Z(n6621) );
  HS65_LS_NAND4ABX3 U16402 ( .A(n5027), .B(n5028), .C(n5029), .D(n5030), .Z(
        n4552) );
  HS65_LS_NOR3X1 U16403 ( .A(n5035), .B(n5036), .C(n5037), .Z(n5029) );
  HS65_LS_NOR4ABX2 U16404 ( .A(n5031), .B(n5032), .C(n5033), .D(n5034), .Z(
        n5030) );
  HS65_LS_OAI212X3 U16405 ( .A(n5038), .B(n5039), .C(n4677), .D(n4488), .E(
        n5040), .Z(n5028) );
  HS65_LS_NAND4ABX3 U16406 ( .A(n8419), .B(n8420), .C(n8421), .D(n8422), .Z(
        n7972) );
  HS65_LS_NOR3X1 U16407 ( .A(n8423), .B(n7803), .C(n8424), .Z(n8422) );
  HS65_LS_OAI222X2 U16408 ( .A(n7833), .B(n7642), .C(n7846), .D(n7687), .E(
        n7818), .F(n8164), .Z(n8420) );
  HS65_LS_NOR3AX2 U16409 ( .A(n8425), .B(n8426), .C(n8427), .Z(n8421) );
  HS65_LS_NAND4ABX3 U16410 ( .A(n8479), .B(n8480), .C(n8481), .D(n8482), .Z(
        n7985) );
  HS65_LS_NOR3X1 U16411 ( .A(n8483), .B(n7903), .C(n8484), .Z(n8482) );
  HS65_LS_OAI222X2 U16412 ( .A(n7932), .B(n7670), .C(n7885), .D(n7725), .E(
        n7917), .F(n8196), .Z(n8480) );
  HS65_LS_NOR3AX2 U16413 ( .A(n8485), .B(n8486), .C(n8487), .Z(n8481) );
  HS65_LS_NOR2X2 U16414 ( .A(n6528), .B(n6337), .Z(n6936) );
  HS65_LS_NOR2X2 U16415 ( .A(n4935), .B(n4744), .Z(n5344) );
  HS65_LS_NOR2X2 U16416 ( .A(n4989), .B(n4783), .Z(n5459) );
  HS65_LS_NOR2X2 U16417 ( .A(n6582), .B(n6376), .Z(n7051) );
  HS65_LS_NOR2X2 U16418 ( .A(n6452), .B(n6230), .Z(n6820) );
  HS65_LS_NOR2X2 U16419 ( .A(n4859), .B(n4637), .Z(n5228) );
  HS65_LS_NAND4ABX3 U16420 ( .A(n3831), .B(n3832), .C(n3833), .D(n3834), .Z(
        n3180) );
  HS65_LS_NOR3X1 U16421 ( .A(n3839), .B(n3840), .C(n3841), .Z(n3833) );
  HS65_LS_OAI212X3 U16422 ( .A(n3842), .B(n3843), .C(n3005), .D(n2848), .E(
        n3844), .Z(n3832) );
  HS65_LS_NOR4ABX2 U16423 ( .A(n3835), .B(n3836), .C(n3837), .D(n3838), .Z(
        n3834) );
  HS65_LS_NOR2X2 U16424 ( .A(n6313), .B(n6152), .Z(n6715) );
  HS65_LS_NOR2X2 U16425 ( .A(n4720), .B(n4559), .Z(n5122) );
  HS65_LS_NAND2X2 U16426 ( .A(n6184), .B(n73), .Z(n6344) );
  HS65_LS_NAND2X2 U16427 ( .A(n4616), .B(n471), .Z(n4790) );
  HS65_LS_NAND2X2 U16428 ( .A(n6209), .B(n294), .Z(n6383) );
  HS65_LS_NAND2X2 U16429 ( .A(n4591), .B(n252), .Z(n4751) );
  HS65_LS_NAND2X2 U16430 ( .A(n4531), .B(n711), .Z(n4644) );
  HS65_LS_NAND2X2 U16431 ( .A(n6124), .B(n529), .Z(n6237) );
  HS65_LS_NOR2X2 U16432 ( .A(n1128), .B(n1399), .Z(n1274) );
  HS65_LS_NAND2X2 U16433 ( .A(n6188), .B(n6057), .Z(n6922) );
  HS65_LS_NAND2X2 U16434 ( .A(n4595), .B(n4464), .Z(n5330) );
  HS65_LS_NAND2X2 U16435 ( .A(n4620), .B(n4510), .Z(n5445) );
  HS65_LS_NAND2X2 U16436 ( .A(n6213), .B(n6103), .Z(n7037) );
  HS65_LS_NAND2X2 U16437 ( .A(n6619), .B(n6081), .Z(n6685) );
  HS65_LS_NAND2X2 U16438 ( .A(n6740), .B(n6137), .Z(n6806) );
  HS65_LS_NAND2X2 U16439 ( .A(n5026), .B(n4488), .Z(n5092) );
  HS65_LS_NAND2X2 U16440 ( .A(n5148), .B(n4544), .Z(n5214) );
  HS65_LS_NOR2X2 U16441 ( .A(n7858), .B(n8663), .Z(n8006) );
  HS65_LS_IVX2 U16442 ( .A(n3101), .Z(n201) );
  HS65_LS_NOR2X2 U16443 ( .A(n7861), .B(n8663), .Z(n8133) );
  HS65_LS_IVX2 U16444 ( .A(n3208), .Z(n420) );
  HS65_LS_NAND2X2 U16445 ( .A(n3002), .B(n3391), .Z(n3828) );
  HS65_LS_NAND2X2 U16446 ( .A(n3454), .B(n3101), .Z(n3468) );
  HS65_LS_NAND2X2 U16447 ( .A(n2984), .B(n3329), .Z(n3711) );
  HS65_LS_NOR2X2 U16448 ( .A(n1880), .B(n2151), .Z(n2026) );
  HS65_LS_NOR3X1 U16449 ( .A(n1819), .B(n1501), .C(n1763), .Z(n1816) );
  HS65_LS_OAI21X2 U16450 ( .A(n1576), .B(n1549), .C(n1771), .Z(n1819) );
  HS65_LS_NOR3X1 U16451 ( .A(n2571), .B(n2253), .C(n2515), .Z(n2568) );
  HS65_LS_OAI21X2 U16452 ( .A(n2328), .B(n2301), .C(n2523), .Z(n2571) );
  HS65_LS_NOR2X2 U16453 ( .A(n8379), .B(n8571), .Z(n8591) );
  HS65_LS_IVX2 U16454 ( .A(n3057), .Z(n152) );
  HS65_LS_NOR2X2 U16455 ( .A(n8315), .B(n8267), .Z(n8222) );
  HS65_LS_NOR2X2 U16456 ( .A(n3146), .B(n3778), .Z(n3336) );
  HS65_LS_NOR2X2 U16457 ( .A(n6080), .B(n6154), .Z(n6675) );
  HS65_LS_NOR2X2 U16458 ( .A(n4487), .B(n4561), .Z(n5082) );
  HS65_LS_NAND4ABX3 U16459 ( .A(n6516), .B(n6517), .C(n6518), .D(n6519), .Z(
        n6189) );
  HS65_LS_OAI222X2 U16460 ( .A(n6528), .B(n6059), .C(n6529), .D(n6338), .E(
        n6056), .F(n6051), .Z(n6517) );
  HS65_LS_NOR4ABX2 U16461 ( .A(n6524), .B(n6525), .C(n6526), .D(n6527), .Z(
        n6518) );
  HS65_LS_NOR4ABX2 U16462 ( .A(n6520), .B(n6521), .C(n6522), .D(n6523), .Z(
        n6519) );
  HS65_LS_NAND4ABX3 U16463 ( .A(n6570), .B(n6571), .C(n6572), .D(n6573), .Z(
        n6201) );
  HS65_LS_OAI222X2 U16464 ( .A(n6582), .B(n6105), .C(n6583), .D(n6377), .E(
        n6102), .F(n6097), .Z(n6571) );
  HS65_LS_NOR4ABX2 U16465 ( .A(n6578), .B(n6579), .C(n6580), .D(n6581), .Z(
        n6572) );
  HS65_LS_NOR4ABX2 U16466 ( .A(n6574), .B(n6575), .C(n6576), .D(n6577), .Z(
        n6573) );
  HS65_LS_NAND4ABX3 U16467 ( .A(n4977), .B(n4978), .C(n4979), .D(n4980), .Z(
        n4608) );
  HS65_LS_OAI222X2 U16468 ( .A(n4989), .B(n4512), .C(n4990), .D(n4784), .E(
        n4509), .F(n4504), .Z(n4978) );
  HS65_LS_NOR4ABX2 U16469 ( .A(n4985), .B(n4986), .C(n4987), .D(n4988), .Z(
        n4979) );
  HS65_LS_NOR4ABX2 U16470 ( .A(n4981), .B(n4982), .C(n4983), .D(n4984), .Z(
        n4980) );
  HS65_LS_NAND4ABX3 U16471 ( .A(n4923), .B(n4924), .C(n4925), .D(n4926), .Z(
        n4596) );
  HS65_LS_OAI222X2 U16472 ( .A(n4935), .B(n4466), .C(n4936), .D(n4745), .E(
        n4463), .F(n4458), .Z(n4924) );
  HS65_LS_NOR4ABX2 U16473 ( .A(n4931), .B(n4932), .C(n4933), .D(n4934), .Z(
        n4925) );
  HS65_LS_NOR4ABX2 U16474 ( .A(n4927), .B(n4928), .C(n4929), .D(n4930), .Z(
        n4926) );
  HS65_LS_NAND4ABX3 U16475 ( .A(n4847), .B(n4848), .C(n4849), .D(n4850), .Z(
        n4538) );
  HS65_LS_OAI222X2 U16476 ( .A(n4859), .B(n4860), .C(n4861), .D(n4638), .E(
        n4862), .F(n4820), .Z(n4848) );
  HS65_LS_NOR4ABX2 U16477 ( .A(n4855), .B(n4856), .C(n4857), .D(n4858), .Z(
        n4849) );
  HS65_LS_NOR4ABX2 U16478 ( .A(n4851), .B(n4852), .C(n4853), .D(n4854), .Z(
        n4850) );
  HS65_LS_NAND4ABX3 U16479 ( .A(n6440), .B(n6441), .C(n6442), .D(n6443), .Z(
        n6131) );
  HS65_LS_OAI222X2 U16480 ( .A(n6452), .B(n6453), .C(n6454), .D(n6231), .E(
        n6455), .F(n6413), .Z(n6441) );
  HS65_LS_NOR4ABX2 U16481 ( .A(n6448), .B(n6449), .C(n6450), .D(n6451), .Z(
        n6442) );
  HS65_LS_NOR4ABX2 U16482 ( .A(n6444), .B(n6445), .C(n6446), .D(n6447), .Z(
        n6443) );
  HS65_LS_NAND4ABX3 U16483 ( .A(n4707), .B(n4708), .C(n4709), .D(n4710), .Z(
        n4482) );
  HS65_LS_OAI222X2 U16484 ( .A(n4719), .B(n4720), .C(n4721), .D(n4561), .E(
        n4680), .F(n4722), .Z(n4708) );
  HS65_LS_NOR4ABX2 U16485 ( .A(n4715), .B(n4716), .C(n4717), .D(n4718), .Z(
        n4709) );
  HS65_LS_NOR4ABX2 U16486 ( .A(n4711), .B(n4712), .C(n4713), .D(n4714), .Z(
        n4710) );
  HS65_LS_NAND4ABX3 U16487 ( .A(n6300), .B(n6301), .C(n6302), .D(n6303), .Z(
        n6075) );
  HS65_LS_OAI222X2 U16488 ( .A(n6312), .B(n6313), .C(n6314), .D(n6154), .E(
        n6273), .F(n6315), .Z(n6301) );
  HS65_LS_NOR4ABX2 U16489 ( .A(n6308), .B(n6309), .C(n6310), .D(n6311), .Z(
        n6302) );
  HS65_LS_NOR4ABX2 U16490 ( .A(n6304), .B(n6305), .C(n6306), .D(n6307), .Z(
        n6303) );
  HS65_LS_NOR2X2 U16491 ( .A(n8149), .B(n7642), .Z(n7798) );
  HS65_LS_NOR2X2 U16492 ( .A(n8181), .B(n7670), .Z(n7898) );
  HS65_LS_NOR2X2 U16493 ( .A(n3189), .B(n2841), .Z(n3397) );
  HS65_LS_NOR2X2 U16494 ( .A(n3148), .B(n2886), .Z(n3335) );
  HS65_LS_NAND2X2 U16495 ( .A(n6084), .B(n573), .Z(n6160) );
  HS65_LS_NAND2X2 U16496 ( .A(n4491), .B(n47), .Z(n4567) );
  HS65_LS_NOR2X2 U16497 ( .A(n3893), .B(n3845), .Z(n3816) );
  HS65_LS_NAND2X2 U16498 ( .A(n6184), .B(n88), .Z(n6531) );
  HS65_LS_NAND2X2 U16499 ( .A(n6209), .B(n309), .Z(n6585) );
  HS65_LS_NAND2X2 U16500 ( .A(n4616), .B(n486), .Z(n4992) );
  HS65_LS_NAND2X2 U16501 ( .A(n4591), .B(n267), .Z(n4938) );
  HS65_LS_NAND2X2 U16502 ( .A(n4531), .B(n705), .Z(n4864) );
  HS65_LS_NAND2X2 U16503 ( .A(n6124), .B(n523), .Z(n6457) );
  HS65_LS_NAND2X2 U16504 ( .A(n4491), .B(n41), .Z(n4724) );
  HS65_LS_NAND2X2 U16505 ( .A(n6084), .B(n567), .Z(n6317) );
  HS65_LS_NAND2X2 U16506 ( .A(n7953), .B(n8525), .Z(n7958) );
  HS65_LS_NOR2X2 U16507 ( .A(n6872), .B(n6050), .Z(n6893) );
  HS65_LS_NOR2X2 U16508 ( .A(n5395), .B(n4503), .Z(n5416) );
  HS65_LS_NOR2X2 U16509 ( .A(n6987), .B(n6096), .Z(n7008) );
  HS65_LS_NOR2X2 U16510 ( .A(n5280), .B(n4457), .Z(n5301) );
  HS65_LS_NOR2X2 U16511 ( .A(n5163), .B(n4835), .Z(n5185) );
  HS65_LS_NOR2X2 U16512 ( .A(n6755), .B(n6428), .Z(n6777) );
  HS65_LS_IVX2 U16513 ( .A(n4676), .Z(n23) );
  HS65_LS_IVX2 U16514 ( .A(n6269), .Z(n549) );
  HS65_LS_AOI12X2 U16515 ( .A(n7686), .B(n8699), .C(n7833), .Z(n9060) );
  HS65_LS_AOI12X2 U16516 ( .A(n7724), .B(n8787), .C(n7932), .Z(n9118) );
  HS65_LS_IVX2 U16517 ( .A(n3297), .Z(n153) );
  HS65_LS_NOR2X2 U16518 ( .A(n2301), .B(n2249), .Z(n2377) );
  HS65_LS_NOR2X2 U16519 ( .A(n1549), .B(n1497), .Z(n1625) );
  HS65_LS_IVX2 U16520 ( .A(n2301), .Z(n898) );
  HS65_LS_IVX2 U16521 ( .A(n1549), .Z(n816) );
  HS65_LS_NAND2X2 U16522 ( .A(n6619), .B(n6314), .Z(n6616) );
  HS65_LS_NAND2X2 U16523 ( .A(n5026), .B(n4721), .Z(n5023) );
  HS65_LS_NAND2X2 U16524 ( .A(n6188), .B(n6529), .Z(n6855) );
  HS65_LS_NAND2X2 U16525 ( .A(n4595), .B(n4936), .Z(n5263) );
  HS65_LS_NAND2X2 U16526 ( .A(n4620), .B(n4990), .Z(n5378) );
  HS65_LS_NAND2X2 U16527 ( .A(n6213), .B(n6583), .Z(n6970) );
  HS65_LS_NAND2X2 U16528 ( .A(n5148), .B(n4861), .Z(n5145) );
  HS65_LS_NAND2X2 U16529 ( .A(n6740), .B(n6454), .Z(n6737) );
  HS65_LS_NAND4ABX3 U16530 ( .A(n8403), .B(n8404), .C(n8405), .D(n8406), .Z(
        n7971) );
  HS65_LS_OAI222X2 U16531 ( .A(n8412), .B(n7842), .C(n8150), .D(n8159), .E(
        n7687), .F(n7686), .Z(n8404) );
  HS65_LS_NOR4ABX2 U16532 ( .A(n7835), .B(n8409), .C(n595), .D(n8410), .Z(
        n8405) );
  HS65_LS_NOR4ABX2 U16533 ( .A(n8407), .B(n7698), .C(n7809), .D(n8408), .Z(
        n8406) );
  HS65_LS_NAND4ABX3 U16534 ( .A(n8463), .B(n8464), .C(n8465), .D(n8466), .Z(
        n7984) );
  HS65_LS_OAI222X2 U16535 ( .A(n8472), .B(n7881), .C(n8182), .D(n8191), .E(
        n7725), .F(n7724), .Z(n8464) );
  HS65_LS_NOR4ABX2 U16536 ( .A(n7934), .B(n8469), .C(n108), .D(n8470), .Z(
        n8465) );
  HS65_LS_NOR4ABX2 U16537 ( .A(n8467), .B(n7736), .C(n7909), .D(n8468), .Z(
        n8466) );
  HS65_LS_OAI21X2 U16538 ( .A(n7777), .B(n8379), .C(n8631), .Z(n8630) );
  HS65_LS_NOR2X2 U16539 ( .A(n1173), .B(n1121), .Z(n1249) );
  HS65_LS_NOR2X2 U16540 ( .A(n1925), .B(n1873), .Z(n2001) );
  HS65_LS_NOR2X2 U16541 ( .A(n6194), .B(n6338), .Z(n6912) );
  HS65_LS_NOR2X2 U16542 ( .A(n4601), .B(n4745), .Z(n5320) );
  HS65_LS_NOR2X2 U16543 ( .A(n4613), .B(n4784), .Z(n5435) );
  HS65_LS_NOR2X2 U16544 ( .A(n6206), .B(n6377), .Z(n7027) );
  HS65_LS_NOR2X2 U16545 ( .A(n4543), .B(n4638), .Z(n5204) );
  HS65_LS_NOR2X2 U16546 ( .A(n6136), .B(n6231), .Z(n6796) );
  HS65_LS_AOI212X2 U16547 ( .A(n839), .B(n818), .C(n847), .D(n823), .E(n1496), 
        .Z(n1495) );
  HS65_LS_OAI21X2 U16548 ( .A(n1497), .B(n1498), .C(n1499), .Z(n1496) );
  HS65_LS_AOI212X2 U16549 ( .A(n921), .B(n900), .C(n929), .D(n905), .E(n2248), 
        .Z(n2247) );
  HS65_LS_OAI21X2 U16550 ( .A(n2249), .B(n2250), .C(n2251), .Z(n2248) );
  HS65_LS_IVX2 U16551 ( .A(n1173), .Z(n857) );
  HS65_LS_IVX2 U16552 ( .A(n4561), .Z(n47) );
  HS65_LS_IVX2 U16553 ( .A(n6154), .Z(n573) );
  HS65_LS_NOR2X2 U16554 ( .A(n2946), .B(n2973), .Z(n3108) );
  HS65_LS_IVX2 U16555 ( .A(n3053), .Z(n179) );
  HS65_LS_IVX2 U16556 ( .A(n1925), .Z(n775) );
  HS65_LS_OAI21X2 U16557 ( .A(n2841), .B(n2842), .C(n2843), .Z(n2840) );
  HS65_LS_NOR2X2 U16558 ( .A(n2299), .B(n2262), .Z(n2489) );
  HS65_LS_NOR2X2 U16559 ( .A(n1547), .B(n1510), .Z(n1737) );
  HS65_LS_OAI21X2 U16560 ( .A(n2886), .B(n2887), .C(n2888), .Z(n2885) );
  HS65_LS_NOR2X2 U16561 ( .A(n8019), .B(n7760), .Z(n8125) );
  HS65_LS_NOR2X2 U16562 ( .A(n8061), .B(n7777), .Z(n8367) );
  HS65_LS_NAND2X2 U16563 ( .A(n612), .B(n7709), .Z(n8155) );
  HS65_LS_NAND2X2 U16564 ( .A(n125), .B(n7747), .Z(n8187) );
  HS65_LS_NAND2X2 U16565 ( .A(n558), .B(n6084), .Z(n6624) );
  HS65_LS_NAND2X2 U16566 ( .A(n32), .B(n4491), .Z(n5031) );
  HS65_LS_IVX2 U16567 ( .A(n4784), .Z(n471) );
  HS65_LS_IVX2 U16568 ( .A(n4745), .Z(n252) );
  HS65_LS_IVX2 U16569 ( .A(n4638), .Z(n711) );
  HS65_LS_IVX2 U16570 ( .A(n6377), .Z(n294) );
  HS65_LS_IVX2 U16571 ( .A(n6338), .Z(n73) );
  HS65_LS_IVX2 U16572 ( .A(n6231), .Z(n529) );
  HS65_LS_NOR2X2 U16573 ( .A(n3391), .B(n2849), .Z(n3408) );
  HS65_LS_NOR2X2 U16574 ( .A(n1171), .B(n1134), .Z(n1361) );
  HS65_LS_NOR2X2 U16575 ( .A(n1923), .B(n1886), .Z(n2113) );
  HS65_LS_OAI212X3 U16576 ( .A(n7831), .B(n7634), .C(n7832), .D(n7833), .E(
        n7834), .Z(n7830) );
  HS65_LS_NOR3X1 U16577 ( .A(n606), .B(n612), .C(n611), .Z(n7831) );
  HS65_LS_OAI21X2 U16578 ( .A(n593), .B(n586), .C(n619), .Z(n7834) );
  HS65_LS_NOR2X2 U16579 ( .A(n7998), .B(n7871), .Z(n8210) );
  HS65_LS_OAI212X3 U16580 ( .A(n4126), .B(n3063), .C(n3599), .D(n3280), .E(
        n4127), .Z(n4125) );
  HS65_LS_NOR3X1 U16581 ( .A(n169), .B(n179), .C(n181), .Z(n4126) );
  HS65_LS_OAI21X2 U16582 ( .A(n155), .B(n150), .C(n175), .Z(n4127) );
  HS65_LS_AOI12X2 U16583 ( .A(n181), .B(n2922), .C(n4171), .Z(n4170) );
  HS65_LS_AOI12X2 U16584 ( .A(n3063), .B(n3282), .C(n3236), .Z(n4171) );
  HS65_LS_NOR2X2 U16585 ( .A(n3187), .B(n2854), .Z(n3815) );
  HS65_LS_OAI21X2 U16586 ( .A(n2973), .B(n3123), .C(n4067), .Z(n4178) );
  HS65_LS_AOI12X2 U16587 ( .A(n430), .B(n2852), .C(n2853), .Z(n2851) );
  HS65_LS_AOI12X2 U16588 ( .A(n2854), .B(n2855), .C(n2856), .Z(n2853) );
  HS65_LS_AOI12X2 U16589 ( .A(n390), .B(n7875), .C(n8673), .Z(n8672) );
  HS65_LS_AOI12X2 U16590 ( .A(n8252), .B(n7870), .C(n8080), .Z(n8673) );
  HS65_LS_AOI12X2 U16591 ( .A(n349), .B(n7958), .C(n8641), .Z(n8640) );
  HS65_LS_AOI12X2 U16592 ( .A(n8556), .B(n7953), .C(n8335), .Z(n8641) );
  HS65_LS_NOR2X2 U16593 ( .A(n3329), .B(n2894), .Z(n3346) );
  HS65_LS_NOR2X2 U16594 ( .A(n3101), .B(n3100), .Z(n3119) );
  HS65_LS_NOR2X2 U16595 ( .A(n8018), .B(n8252), .Z(n8221) );
  HS65_LS_NOR2X2 U16596 ( .A(n8060), .B(n8556), .Z(n8526) );
  HS65_LS_NAND2X2 U16597 ( .A(n574), .B(n6084), .Z(n6644) );
  HS65_LS_NAND2X2 U16598 ( .A(n48), .B(n4491), .Z(n5051) );
  HS65_LS_AOI12X2 U16599 ( .A(n46), .B(n4579), .C(n4580), .Z(n4578) );
  HS65_LS_AOI12X2 U16600 ( .A(n4581), .B(n4562), .C(n4582), .Z(n4580) );
  HS65_LS_AOI12X2 U16601 ( .A(n572), .B(n6172), .C(n6173), .Z(n6171) );
  HS65_LS_AOI12X2 U16602 ( .A(n6174), .B(n6155), .C(n6175), .Z(n6173) );
  HS65_LS_AOI12X2 U16603 ( .A(n608), .B(n8162), .C(n8163), .Z(n8161) );
  HS65_LS_AOI12X2 U16604 ( .A(n8164), .B(n7646), .C(n7644), .Z(n8163) );
  HS65_LS_AOI12X2 U16605 ( .A(n121), .B(n8194), .C(n8195), .Z(n8193) );
  HS65_LS_AOI12X2 U16606 ( .A(n8196), .B(n7674), .C(n7672), .Z(n8195) );
  HS65_LS_AOI12X2 U16607 ( .A(n857), .B(n1132), .C(n1133), .Z(n1131) );
  HS65_LS_AOI12X2 U16608 ( .A(n1134), .B(n1135), .C(n1136), .Z(n1133) );
  HS65_LS_AOI12X2 U16609 ( .A(n775), .B(n1884), .C(n1885), .Z(n1883) );
  HS65_LS_AOI12X2 U16610 ( .A(n1886), .B(n1887), .C(n1888), .Z(n1885) );
  HS65_LS_AOI12X2 U16611 ( .A(n816), .B(n1508), .C(n1509), .Z(n1507) );
  HS65_LS_AOI12X2 U16612 ( .A(n1510), .B(n1511), .C(n1512), .Z(n1509) );
  HS65_LS_AOI12X2 U16613 ( .A(n898), .B(n2260), .C(n2261), .Z(n2259) );
  HS65_LS_AOI12X2 U16614 ( .A(n2262), .B(n2263), .C(n2264), .Z(n2261) );
  HS65_LS_AOI12X2 U16615 ( .A(n227), .B(n2872), .C(n4233), .Z(n4232) );
  HS65_LS_AOI12X2 U16616 ( .A(n3470), .B(n3905), .C(n3074), .Z(n4233) );
  HS65_LS_NOR2X2 U16617 ( .A(n1243), .B(n1129), .Z(n1260) );
  HS65_LS_NOR2X2 U16618 ( .A(n1995), .B(n1881), .Z(n2012) );
  HS65_LS_NOR2X2 U16619 ( .A(n1619), .B(n1505), .Z(n1636) );
  HS65_LS_NOR2X2 U16620 ( .A(n2371), .B(n2257), .Z(n2388) );
  HS65_LS_AOI12X2 U16621 ( .A(n654), .B(n2897), .C(n2898), .Z(n2896) );
  HS65_LS_AOI12X2 U16622 ( .A(n2899), .B(n2900), .C(n2901), .Z(n2898) );
  HS65_LS_NOR2X2 U16623 ( .A(n4488), .B(n5524), .Z(n5016) );
  HS65_LS_NOR2X2 U16624 ( .A(n6057), .B(n7136), .Z(n6848) );
  HS65_LS_NOR2X2 U16625 ( .A(n4464), .B(n5544), .Z(n5256) );
  HS65_LS_NOR2X2 U16626 ( .A(n4510), .B(n5565), .Z(n5371) );
  HS65_LS_NOR2X2 U16627 ( .A(n6103), .B(n7157), .Z(n6963) );
  HS65_LS_NOR2X2 U16628 ( .A(n6081), .B(n7116), .Z(n6609) );
  HS65_LS_NOR2X2 U16629 ( .A(n6137), .B(n7181), .Z(n6730) );
  HS65_LS_NOR2X2 U16630 ( .A(n4544), .B(n5589), .Z(n5138) );
  HS65_LS_OAI212X3 U16631 ( .A(n2322), .B(n2323), .C(n2324), .D(n2256), .E(
        n2325), .Z(n2318) );
  HS65_LS_AOI12X2 U16632 ( .A(n894), .B(n2326), .C(n2327), .Z(n2325) );
  HS65_LS_AOI12X2 U16633 ( .A(n2328), .B(n2300), .C(n2329), .Z(n2327) );
  HS65_LS_OAI212X3 U16634 ( .A(n1570), .B(n1571), .C(n1572), .D(n1504), .E(
        n1573), .Z(n1566) );
  HS65_LS_AOI12X2 U16635 ( .A(n812), .B(n1574), .C(n1575), .Z(n1573) );
  HS65_LS_AOI12X2 U16636 ( .A(n1576), .B(n1548), .C(n1577), .Z(n1575) );
  HS65_LS_NOR4ABX2 U16637 ( .A(n3906), .B(n3907), .C(n3908), .D(n3909), .Z(
        n3901) );
  HS65_LS_OAI212X3 U16638 ( .A(n3127), .B(n3538), .C(n2946), .D(n2943), .E(
        n3910), .Z(n3909) );
  HS65_LS_AOI12X2 U16639 ( .A(n47), .B(n4497), .C(n5764), .Z(n5763) );
  HS65_LS_AOI12X2 U16640 ( .A(n4495), .B(n5492), .C(n4493), .Z(n5764) );
  HS65_LS_AOI12X2 U16641 ( .A(n573), .B(n6090), .C(n7356), .Z(n7355) );
  HS65_LS_AOI12X2 U16642 ( .A(n6088), .B(n7084), .C(n6086), .Z(n7356) );
  HS65_LS_NAND3X2 U16643 ( .A(n3214), .B(n3415), .C(n3202), .Z(n4052) );
  HS65_LS_AOI12X2 U16644 ( .A(n471), .B(n4514), .C(n4515), .Z(n4513) );
  HS65_LS_AOI12X2 U16645 ( .A(n4516), .B(n4517), .C(n4518), .Z(n4515) );
  HS65_LS_AOI12X2 U16646 ( .A(n252), .B(n4468), .C(n4469), .Z(n4467) );
  HS65_LS_AOI12X2 U16647 ( .A(n4470), .B(n4471), .C(n4472), .Z(n4469) );
  HS65_LS_AOI12X2 U16648 ( .A(n294), .B(n6107), .C(n6108), .Z(n6106) );
  HS65_LS_AOI12X2 U16649 ( .A(n6109), .B(n6110), .C(n6111), .Z(n6108) );
  HS65_LS_AOI12X2 U16650 ( .A(n711), .B(n4537), .C(n5826), .Z(n5825) );
  HS65_LS_AOI12X2 U16651 ( .A(n4535), .B(n5508), .C(n4533), .Z(n5826) );
  HS65_LS_AOI12X2 U16652 ( .A(n529), .B(n6130), .C(n7418), .Z(n7417) );
  HS65_LS_AOI12X2 U16653 ( .A(n6128), .B(n7100), .C(n6126), .Z(n7418) );
  HS65_LS_AOI12X2 U16654 ( .A(n73), .B(n6061), .C(n6062), .Z(n6060) );
  HS65_LS_AOI12X2 U16655 ( .A(n6063), .B(n6064), .C(n6065), .Z(n6062) );
  HS65_LS_AOI12X2 U16656 ( .A(n656), .B(n3165), .C(n3166), .Z(n3164) );
  HS65_LS_AOI12X2 U16657 ( .A(n3167), .B(n3147), .C(n3168), .Z(n3166) );
  HS65_LS_AOI12X2 U16658 ( .A(n474), .B(n4802), .C(n4803), .Z(n4801) );
  HS65_LS_AOI12X2 U16659 ( .A(n4804), .B(n4785), .C(n4805), .Z(n4803) );
  HS65_LS_AOI12X2 U16660 ( .A(n297), .B(n6395), .C(n6396), .Z(n6394) );
  HS65_LS_AOI12X2 U16661 ( .A(n6397), .B(n6378), .C(n6398), .Z(n6396) );
  HS65_LS_NOR2X2 U16662 ( .A(n3146), .B(n2899), .Z(n3698) );
  HS65_LS_NAND3X2 U16663 ( .A(n2971), .B(n3127), .C(n2959), .Z(n3943) );
  HS65_LS_NOR2X2 U16664 ( .A(n6063), .B(n6337), .Z(n6924) );
  HS65_LS_NOR2X2 U16665 ( .A(n4470), .B(n4744), .Z(n5332) );
  HS65_LS_NOR2X2 U16666 ( .A(n4516), .B(n4783), .Z(n5447) );
  HS65_LS_NOR2X2 U16667 ( .A(n6109), .B(n6376), .Z(n7039) );
  HS65_LS_NOR2X2 U16668 ( .A(n6128), .B(n6230), .Z(n6808) );
  HS65_LS_NOR2X2 U16669 ( .A(n4535), .B(n4637), .Z(n5216) );
  HS65_LS_NOR2X2 U16670 ( .A(n6088), .B(n6152), .Z(n6687) );
  HS65_LS_NOR2X2 U16671 ( .A(n4495), .B(n4559), .Z(n5094) );
  HS65_LS_NOR4ABX2 U16672 ( .A(n8859), .B(n8865), .C(n8633), .D(n8888), .Z(
        n8884) );
  HS65_LS_OAI212X3 U16673 ( .A(n8051), .B(n7955), .C(n8556), .D(n8542), .E(
        n7781), .Z(n8888) );
  HS65_LS_AOI12X2 U16674 ( .A(n432), .B(n3206), .C(n3207), .Z(n3205) );
  HS65_LS_AOI12X2 U16675 ( .A(n3208), .B(n3188), .C(n3209), .Z(n3207) );
  HS65_LS_NOR2X2 U16676 ( .A(n3297), .B(n3044), .Z(n3047) );
  HS65_LS_NAND3X2 U16677 ( .A(n7871), .B(n8130), .C(n7997), .Z(n9003) );
  HS65_LS_NAND3X2 U16678 ( .A(n7954), .B(n8326), .C(n8039), .Z(n8943) );
  HS65_LS_NOR2X2 U16679 ( .A(n4680), .B(n4561), .Z(n4728) );
  HS65_LS_NOR2X2 U16680 ( .A(n6273), .B(n6154), .Z(n6321) );
  HS65_LS_NOR2X2 U16681 ( .A(n7724), .B(n8181), .Z(n7923) );
  HS65_LS_NOR2X2 U16682 ( .A(n7686), .B(n8149), .Z(n7824) );
  HS65_LS_NOR2X2 U16683 ( .A(n8186), .B(n8181), .Z(n7919) );
  HS65_LS_NOR2X2 U16684 ( .A(n8154), .B(n8149), .Z(n7820) );
  HS65_LS_AOI12X2 U16685 ( .A(n124), .B(n7883), .C(n7884), .Z(n7882) );
  HS65_LS_AOI12X2 U16686 ( .A(n7662), .B(n7885), .C(n7886), .Z(n7884) );
  HS65_LS_AOI12X2 U16687 ( .A(n611), .B(n7844), .C(n7845), .Z(n7843) );
  HS65_LS_AOI12X2 U16688 ( .A(n7634), .B(n7846), .C(n7847), .Z(n7845) );
  HS65_LS_IVX2 U16689 ( .A(n7959), .Z(n318) );
  HS65_LS_IVX2 U16690 ( .A(n7953), .Z(n334) );
  HS65_LS_NAND2X2 U16691 ( .A(n619), .B(n7709), .Z(n8409) );
  HS65_LS_NAND2X2 U16692 ( .A(n132), .B(n7747), .Z(n8469) );
  HS65_LS_NOR4ABX2 U16693 ( .A(n7865), .B(n7866), .C(n7867), .D(n7868), .Z(
        n7854) );
  HS65_LS_OA212X4 U16694 ( .A(n7869), .B(n7870), .C(n7871), .D(n7872), .E(
        n7873), .Z(n7865) );
  HS65_LS_NOR2X2 U16695 ( .A(n6051), .B(n6338), .Z(n6535) );
  HS65_LS_NOR2X2 U16696 ( .A(n6097), .B(n6377), .Z(n6589) );
  HS65_LS_NOR2X2 U16697 ( .A(n4504), .B(n4784), .Z(n4996) );
  HS65_LS_NOR2X2 U16698 ( .A(n4458), .B(n4745), .Z(n4942) );
  HS65_LS_NOR2X2 U16699 ( .A(n4820), .B(n4638), .Z(n4868) );
  HS65_LS_NOR2X2 U16700 ( .A(n6413), .B(n6231), .Z(n6461) );
  HS65_LS_OAI212X3 U16701 ( .A(n6504), .B(n6050), .C(n6065), .D(n6353), .E(
        n6505), .Z(n6493) );
  HS65_LS_NOR2X2 U16702 ( .A(n56), .B(n55), .Z(n6504) );
  HS65_LS_OAI21X2 U16703 ( .A(n61), .B(n68), .C(n83), .Z(n6505) );
  HS65_LS_OAI212X3 U16704 ( .A(n6558), .B(n6096), .C(n6111), .D(n6392), .E(
        n6559), .Z(n6547) );
  HS65_LS_NOR2X2 U16705 ( .A(n277), .B(n276), .Z(n6558) );
  HS65_LS_OAI21X2 U16706 ( .A(n282), .B(n289), .C(n304), .Z(n6559) );
  HS65_LS_OAI212X3 U16707 ( .A(n4911), .B(n4457), .C(n4472), .D(n4760), .E(
        n4912), .Z(n4900) );
  HS65_LS_NOR2X2 U16708 ( .A(n235), .B(n234), .Z(n4911) );
  HS65_LS_OAI21X2 U16709 ( .A(n240), .B(n247), .C(n262), .Z(n4912) );
  HS65_LS_OAI212X3 U16710 ( .A(n4965), .B(n4503), .C(n4518), .D(n4799), .E(
        n4966), .Z(n4954) );
  HS65_LS_NOR2X2 U16711 ( .A(n454), .B(n453), .Z(n4965) );
  HS65_LS_OAI21X2 U16712 ( .A(n459), .B(n466), .C(n481), .Z(n4966) );
  HS65_LS_OAI212X3 U16713 ( .A(n4834), .B(n4835), .C(n4533), .D(n4653), .E(
        n4836), .Z(n4823) );
  HS65_LS_NOR2X2 U16714 ( .A(n688), .B(n687), .Z(n4834) );
  HS65_LS_OAI21X2 U16715 ( .A(n685), .B(n675), .C(n700), .Z(n4836) );
  HS65_LS_OAI212X3 U16716 ( .A(n6427), .B(n6428), .C(n6126), .D(n6246), .E(
        n6429), .Z(n6416) );
  HS65_LS_NOR2X2 U16717 ( .A(n506), .B(n505), .Z(n6427) );
  HS65_LS_OAI21X2 U16718 ( .A(n503), .B(n493), .C(n518), .Z(n6429) );
  HS65_LS_OAI212X3 U16719 ( .A(n4694), .B(n4695), .C(n4493), .D(n4576), .E(
        n4696), .Z(n4683) );
  HS65_LS_NOR2X2 U16720 ( .A(n24), .B(n23), .Z(n4694) );
  HS65_LS_OAI21X2 U16721 ( .A(n21), .B(n10), .C(n36), .Z(n4696) );
  HS65_LS_OAI212X3 U16722 ( .A(n6287), .B(n6288), .C(n6086), .D(n6169), .E(
        n6289), .Z(n6276) );
  HS65_LS_NOR2X2 U16723 ( .A(n550), .B(n549), .Z(n6287) );
  HS65_LS_OAI21X2 U16724 ( .A(n547), .B(n536), .C(n562), .Z(n6289) );
  HS65_LS_NOR4ABX2 U16725 ( .A(n9024), .B(n8721), .C(n8399), .D(n8757), .Z(
        n9021) );
  HS65_LS_OAI21X2 U16726 ( .A(n584), .B(n7709), .C(n624), .Z(n9024) );
  HS65_LS_NOR4ABX2 U16727 ( .A(n9082), .B(n8809), .C(n8459), .D(n8845), .Z(
        n9079) );
  HS65_LS_OAI21X2 U16728 ( .A(n97), .B(n7747), .C(n137), .Z(n9082) );
  HS65_LS_NOR4ABX2 U16729 ( .A(n5747), .B(n5111), .C(n5080), .D(n4703), .Z(
        n5744) );
  HS65_LS_OAI21X2 U16730 ( .A(n15), .B(n4491), .C(n31), .Z(n5747) );
  HS65_LS_NOR4ABX2 U16731 ( .A(n7339), .B(n6704), .C(n6673), .D(n6296), .Z(
        n7336) );
  HS65_LS_OAI21X2 U16732 ( .A(n541), .B(n6084), .C(n557), .Z(n7339) );
  HS65_LS_NAND4ABX3 U16733 ( .A(n2277), .B(n2293), .C(n2343), .D(n2344), .Z(
        n2331) );
  HS65_LS_AOI212X2 U16734 ( .A(n915), .B(n2345), .C(n908), .D(n916), .E(n2346), 
        .Z(n2344) );
  HS65_LS_OAI21X2 U16735 ( .A(n2249), .B(n2264), .C(n2347), .Z(n2346) );
  HS65_LS_NAND4ABX3 U16736 ( .A(n1525), .B(n1541), .C(n1591), .D(n1592), .Z(
        n1579) );
  HS65_LS_AOI212X2 U16737 ( .A(n833), .B(n1593), .C(n826), .D(n834), .E(n1594), 
        .Z(n1592) );
  HS65_LS_OAI21X2 U16738 ( .A(n1497), .B(n1512), .C(n1595), .Z(n1594) );
  HS65_LS_NAND4ABX3 U16739 ( .A(n1149), .B(n1165), .C(n1215), .D(n1216), .Z(
        n1203) );
  HS65_LS_AOI212X2 U16740 ( .A(n874), .B(n1217), .C(n867), .D(n875), .E(n1218), 
        .Z(n1216) );
  HS65_LS_OAI21X2 U16741 ( .A(n1121), .B(n1136), .C(n1219), .Z(n1218) );
  HS65_LS_NAND4ABX3 U16742 ( .A(n1901), .B(n1917), .C(n1967), .D(n1968), .Z(
        n1955) );
  HS65_LS_AOI212X2 U16743 ( .A(n792), .B(n1969), .C(n785), .D(n793), .E(n1970), 
        .Z(n1968) );
  HS65_LS_OAI21X2 U16744 ( .A(n1873), .B(n1888), .C(n1971), .Z(n1970) );
  HS65_LS_AOI12X2 U16745 ( .A(n1158), .B(n1214), .C(n1156), .Z(n1210) );
  HS65_LS_AOI12X2 U16746 ( .A(n2286), .B(n2342), .C(n2284), .Z(n2338) );
  HS65_LS_AOI12X2 U16747 ( .A(n1910), .B(n1966), .C(n1908), .Z(n1962) );
  HS65_LS_AOI12X2 U16748 ( .A(n1534), .B(n1590), .C(n1532), .Z(n1586) );
  HS65_LS_NOR4ABX2 U16749 ( .A(n5908), .B(n5431), .C(n4973), .D(n5478), .Z(
        n5905) );
  HS65_LS_OAI21X2 U16750 ( .A(n464), .B(n4616), .C(n480), .Z(n5908) );
  HS65_LS_NOR4ABX2 U16751 ( .A(n5849), .B(n5316), .C(n4919), .D(n5363), .Z(
        n5846) );
  HS65_LS_OAI21X2 U16752 ( .A(n245), .B(n4591), .C(n261), .Z(n5849) );
  HS65_LS_NOR4ABX2 U16753 ( .A(n7500), .B(n7023), .C(n6566), .D(n7070), .Z(
        n7497) );
  HS65_LS_OAI21X2 U16754 ( .A(n287), .B(n6209), .C(n303), .Z(n7500) );
  HS65_LS_NOR4ABX2 U16755 ( .A(n5809), .B(n5200), .C(n4843), .D(n5248), .Z(
        n5806) );
  HS65_LS_OAI21X2 U16756 ( .A(n680), .B(n4531), .C(n695), .Z(n5809) );
  HS65_LS_NOR4ABX2 U16757 ( .A(n7401), .B(n6792), .C(n6436), .D(n6840), .Z(
        n7398) );
  HS65_LS_OAI21X2 U16758 ( .A(n498), .B(n6124), .C(n513), .Z(n7401) );
  HS65_LS_NOR4ABX2 U16759 ( .A(n7441), .B(n6908), .C(n6512), .D(n6955), .Z(
        n7438) );
  HS65_LS_OAI21X2 U16760 ( .A(n66), .B(n6184), .C(n82), .Z(n7441) );
  HS65_LS_AOI12X2 U16761 ( .A(n2989), .B(n3359), .C(n2987), .Z(n3355) );
  HS65_LS_AOI12X2 U16762 ( .A(n3007), .B(n3421), .C(n3005), .Z(n3417) );
  HS65_LS_OAI21X2 U16763 ( .A(n6269), .B(n6312), .C(n6699), .Z(n7328) );
  HS65_LS_OAI21X2 U16764 ( .A(n4676), .B(n4719), .C(n5106), .Z(n5736) );
  HS65_LS_OAI21X2 U16765 ( .A(n6487), .B(n6059), .C(n6949), .Z(n7462) );
  HS65_LS_OAI21X2 U16766 ( .A(n5008), .B(n4512), .C(n5472), .Z(n5929) );
  HS65_LS_OAI21X2 U16767 ( .A(n6601), .B(n6105), .C(n7064), .Z(n7521) );
  HS65_LS_OAI21X2 U16768 ( .A(n4894), .B(n4466), .C(n5357), .Z(n5870) );
  HS65_LS_OAI21X2 U16769 ( .A(n4880), .B(n4860), .C(n5242), .Z(n5798) );
  HS65_LS_OAI21X2 U16770 ( .A(n6473), .B(n6453), .C(n6834), .Z(n7390) );
  HS65_LS_NAND2X2 U16771 ( .A(n74), .B(n6184), .Z(n6881) );
  HS65_LS_NAND2X2 U16772 ( .A(n472), .B(n4616), .Z(n5404) );
  HS65_LS_NAND2X2 U16773 ( .A(n712), .B(n4531), .Z(n5172) );
  HS65_LS_NAND2X2 U16774 ( .A(n295), .B(n6209), .Z(n6996) );
  HS65_LS_NAND2X2 U16775 ( .A(n253), .B(n4591), .Z(n5289) );
  HS65_LS_NAND2X2 U16776 ( .A(n530), .B(n6124), .Z(n6764) );
  HS65_LS_NAND2X2 U16777 ( .A(n609), .B(n7709), .Z(n7706) );
  HS65_LS_NAND2X2 U16778 ( .A(n122), .B(n7747), .Z(n7744) );
  HS65_LS_NAND2X2 U16779 ( .A(n6194), .B(n6529), .Z(n6940) );
  HS65_LS_NAND2X2 U16780 ( .A(n4601), .B(n4936), .Z(n5348) );
  HS65_LS_NAND2X2 U16781 ( .A(n4613), .B(n4990), .Z(n5463) );
  HS65_LS_NAND2X2 U16782 ( .A(n6206), .B(n6583), .Z(n7055) );
  HS65_LS_NAND2X2 U16783 ( .A(n6136), .B(n6454), .Z(n6824) );
  HS65_LS_NAND2X2 U16784 ( .A(n4543), .B(n4861), .Z(n5232) );
  HS65_LS_NAND2X2 U16785 ( .A(n8525), .B(n7964), .Z(n8523) );
  HS65_LS_OAI21X2 U16786 ( .A(n8154), .B(n7842), .C(n8759), .Z(n9019) );
  HS65_LS_OAI21X2 U16787 ( .A(n8186), .B(n7881), .C(n8847), .Z(n9077) );
  HS65_LS_NAND2X2 U16788 ( .A(n7747), .B(n135), .Z(n7934) );
  HS65_LS_NAND2X2 U16789 ( .A(n7709), .B(n622), .Z(n7835) );
  HS65_LS_NAND2X2 U16790 ( .A(n8525), .B(n8069), .Z(n8554) );
  HS65_LS_NAND2X2 U16791 ( .A(n4616), .B(n478), .Z(n4985) );
  HS65_LS_NAND2X2 U16792 ( .A(n4591), .B(n259), .Z(n4931) );
  HS65_LS_NAND2X2 U16793 ( .A(n6209), .B(n301), .Z(n6578) );
  HS65_LS_NAND2X2 U16794 ( .A(n4531), .B(n697), .Z(n4855) );
  HS65_LS_NAND2X2 U16795 ( .A(n6124), .B(n515), .Z(n6448) );
  HS65_LS_NAND2X2 U16796 ( .A(n6184), .B(n80), .Z(n6524) );
  HS65_LS_NAND2X2 U16797 ( .A(n4491), .B(n33), .Z(n4715) );
  HS65_LS_NAND2X2 U16798 ( .A(n6084), .B(n559), .Z(n6308) );
  HS65_LS_NAND2X2 U16799 ( .A(n6080), .B(n6314), .Z(n6719) );
  HS65_LS_NAND2X2 U16800 ( .A(n4487), .B(n4721), .Z(n5126) );
  HS65_LS_NAND2X2 U16801 ( .A(n7735), .B(n8191), .Z(n8839) );
  HS65_LS_NAND2X2 U16802 ( .A(n7697), .B(n8159), .Z(n8751) );
  HS65_LS_AOI12X2 U16803 ( .A(n43), .B(n4671), .C(n5653), .Z(n5652) );
  HS65_LS_AOI12X2 U16804 ( .A(n4680), .B(n5526), .C(n4722), .Z(n5653) );
  HS65_LS_AOI12X2 U16805 ( .A(n569), .B(n6264), .C(n7245), .Z(n7244) );
  HS65_LS_AOI12X2 U16806 ( .A(n6273), .B(n7118), .C(n6315), .Z(n7245) );
  HS65_LS_AOI12X2 U16807 ( .A(n358), .B(n7775), .C(n7776), .Z(n7772) );
  HS65_LS_AOI12X2 U16808 ( .A(n7777), .B(n7778), .C(n7779), .Z(n7776) );
  HS65_LS_AOI12X2 U16809 ( .A(n620), .B(n7684), .C(n7685), .Z(n7681) );
  HS65_LS_AOI12X2 U16810 ( .A(n7686), .B(n7642), .C(n7687), .Z(n7685) );
  HS65_LS_AOI12X2 U16811 ( .A(n133), .B(n7722), .C(n7723), .Z(n7719) );
  HS65_LS_AOI12X2 U16812 ( .A(n7724), .B(n7670), .C(n7725), .Z(n7723) );
  HS65_LS_AOI12X2 U16813 ( .A(n395), .B(n7758), .C(n7759), .Z(n7755) );
  HS65_LS_AOI12X2 U16814 ( .A(n7760), .B(n7761), .C(n7762), .Z(n7759) );
  HS65_LS_OAI212X3 U16815 ( .A(n3894), .B(n2841), .C(n3005), .D(n3391), .E(
        n4051), .Z(n4049) );
  HS65_LS_CB4I1X4 U16816 ( .A(n3985), .B(n3215), .C(n3845), .D(n3896), .Z(
        n4051) );
  HS65_LS_CB4I1X4 U16817 ( .A(n1780), .B(n1777), .C(n1688), .D(n1754), .Z(
        n1804) );
  HS65_LS_CB4I1X4 U16818 ( .A(n2532), .B(n2529), .C(n2440), .D(n2506), .Z(
        n2556) );
  HS65_LS_CB4I1X4 U16819 ( .A(n1404), .B(n1401), .C(n1312), .D(n1378), .Z(
        n1428) );
  HS65_LS_CB4I1X4 U16820 ( .A(n3942), .B(n2972), .C(n3486), .D(n3539), .Z(
        n3941) );
  HS65_LS_CB4I1X4 U16821 ( .A(n2156), .B(n2153), .C(n2064), .D(n2130), .Z(
        n2180) );
  HS65_LS_CB4I1X4 U16822 ( .A(n3964), .B(n3174), .C(n3728), .D(n3779), .Z(
        n4027) );
  HS65_LS_CB4I1X4 U16823 ( .A(n8881), .B(n8051), .C(n8571), .D(n8544), .Z(
        n8937) );
  HS65_LS_MX41X4 U16824 ( .D0(n551), .S0(n574), .D1(n547), .S1(n557), .D2(n564), .S2(n6084), .D3(n569), .S3(n549), .Z(n6680) );
  HS65_LS_MX41X4 U16825 ( .D0(n25), .S0(n48), .D1(n21), .S1(n31), .D2(n38), 
        .S2(n4491), .D3(n43), .S3(n23), .Z(n5087) );
  HS65_LS_MX41X4 U16826 ( .D0(n106), .S0(n122), .D1(n137), .S1(n114), .D2(n126), .S2(n7747), .D3(n110), .S3(n133), .Z(n8820) );
  HS65_LS_MX41X4 U16827 ( .D0(n593), .S0(n609), .D1(n624), .S1(n601), .D2(n613), .S2(n7709), .D3(n597), .S3(n620), .Z(n8732) );
  HS65_LS_MX41X4 U16828 ( .D0(n57), .S0(n74), .D1(n61), .S1(n82), .D2(n84), 
        .S2(n6184), .D3(n87), .S3(n55), .Z(n6917) );
  HS65_LS_MX41X4 U16829 ( .D0(n236), .S0(n253), .D1(n240), .S1(n261), .D2(n263), .S2(n4591), .D3(n266), .S3(n234), .Z(n5325) );
  HS65_LS_MX41X4 U16830 ( .D0(n455), .S0(n472), .D1(n459), .S1(n480), .D2(n482), .S2(n4616), .D3(n485), .S3(n453), .Z(n5440) );
  HS65_LS_MX41X4 U16831 ( .D0(n278), .S0(n295), .D1(n282), .S1(n303), .D2(n305), .S2(n6209), .D3(n308), .S3(n276), .Z(n7032) );
  HS65_LS_MX41X4 U16832 ( .D0(n507), .S0(n530), .D1(n503), .S1(n513), .D2(n520), .S2(n6124), .D3(n525), .S3(n505), .Z(n6801) );
  HS65_LS_MX41X4 U16833 ( .D0(n689), .S0(n712), .D1(n685), .S1(n695), .D2(n702), .S2(n4531), .D3(n707), .S3(n687), .Z(n5209) );
  HS65_LS_OA12X4 U16834 ( .A(n8525), .B(n7961), .C(n8601), .Z(n8600) );
  HS65_LS_NAND2X2 U16835 ( .A(n3067), .B(n2927), .Z(n3292) );
  HS65_LS_AOI12X2 U16836 ( .A(n7777), .B(n8571), .C(n8070), .Z(n8880) );
  HS65_LS_AOI12X2 U16837 ( .A(n3067), .B(n3625), .C(n3280), .Z(n3922) );
  HS65_LS_OAI21X2 U16838 ( .A(n3536), .B(n3126), .C(n4059), .Z(n4058) );
  HS65_LS_OAI21X2 U16839 ( .A(n191), .B(n193), .C(n219), .Z(n4059) );
  HS65_LS_AOI12X2 U16840 ( .A(n7760), .B(n8267), .C(n8031), .Z(n8507) );
  HS65_LS_AOI12X2 U16841 ( .A(n6413), .B(n6755), .C(n6753), .Z(n7098) );
  HS65_LS_AOI12X2 U16842 ( .A(n4680), .B(n5041), .C(n5039), .Z(n5490) );
  HS65_LS_AOI12X2 U16843 ( .A(n6273), .B(n6634), .C(n6632), .Z(n7082) );
  HS65_LS_AOI12X2 U16844 ( .A(n4820), .B(n5163), .C(n5161), .Z(n5506) );
  HS65_LS_AOI12X2 U16845 ( .A(n4533), .B(n4534), .C(n4535), .Z(n4532) );
  HS65_LS_AOI12X2 U16846 ( .A(n4518), .B(n4618), .C(n4516), .Z(n4617) );
  HS65_LS_AOI12X2 U16847 ( .A(n6111), .B(n6211), .C(n6109), .Z(n6210) );
  HS65_LS_AOI12X2 U16848 ( .A(n6065), .B(n6186), .C(n6063), .Z(n6185) );
  HS65_LS_AOI12X2 U16849 ( .A(n6126), .B(n6127), .C(n6128), .Z(n6125) );
  HS65_LS_AOI12X2 U16850 ( .A(n4472), .B(n4593), .C(n4470), .Z(n4592) );
  HS65_LS_AOI12X2 U16851 ( .A(n2973), .B(n3486), .C(n3484), .Z(n3912) );
  HS65_LS_AOI12X2 U16852 ( .A(n7847), .B(n7978), .C(n7634), .Z(n7977) );
  HS65_LS_AOI12X2 U16853 ( .A(n7886), .B(n7991), .C(n7662), .Z(n7990) );
  HS65_LS_AOI12X2 U16854 ( .A(n6086), .B(n6087), .C(n6088), .Z(n6085) );
  HS65_LS_AOI12X2 U16855 ( .A(n4493), .B(n4494), .C(n4495), .Z(n4492) );
  HS65_LS_AOI12X2 U16856 ( .A(n4487), .B(n4676), .C(n4677), .Z(n4672) );
  HS65_LS_AOI12X2 U16857 ( .A(n6080), .B(n6269), .C(n6270), .Z(n6265) );
  HS65_LS_AOI12X2 U16858 ( .A(n4543), .B(n4880), .C(n4881), .Z(n4876) );
  HS65_LS_AOI12X2 U16859 ( .A(n6136), .B(n6473), .C(n6474), .Z(n6469) );
  HS65_LS_NAND2X2 U16860 ( .A(n4680), .B(n4487), .Z(n4671) );
  HS65_LS_NAND2X2 U16861 ( .A(n6273), .B(n6080), .Z(n6264) );
  HS65_LS_AOI12X2 U16862 ( .A(n3042), .B(n3063), .C(n3064), .Z(n3060) );
  HS65_LS_AOI12X2 U16863 ( .A(n7697), .B(n8154), .C(n8436), .Z(n8432) );
  HS65_LS_AOI12X2 U16864 ( .A(n7735), .B(n8186), .C(n8447), .Z(n8443) );
  HS65_LS_AOI12X2 U16865 ( .A(n2927), .B(n3297), .C(n2925), .Z(n3293) );
  HS65_LS_AOI12X2 U16866 ( .A(n180), .B(n3055), .C(n3056), .Z(n3054) );
  HS65_LS_AOI12X2 U16867 ( .A(n3057), .B(n3045), .C(n3058), .Z(n3056) );
  HS65_LS_AOI12X2 U16868 ( .A(n387), .B(n8001), .C(n8002), .Z(n8000) );
  HS65_LS_AOI12X2 U16869 ( .A(n8003), .B(n8004), .C(n7869), .Z(n8002) );
  HS65_LS_AOI12X2 U16870 ( .A(n76), .B(n6356), .C(n6357), .Z(n6355) );
  HS65_LS_AOI12X2 U16871 ( .A(n6358), .B(n6339), .C(n6359), .Z(n6357) );
  HS65_LS_AOI12X2 U16872 ( .A(n255), .B(n4763), .C(n4764), .Z(n4762) );
  HS65_LS_AOI12X2 U16873 ( .A(n4765), .B(n4746), .C(n4766), .Z(n4764) );
  HS65_LS_AOI12X2 U16874 ( .A(n710), .B(n4656), .C(n4657), .Z(n4655) );
  HS65_LS_AOI12X2 U16875 ( .A(n4658), .B(n4639), .C(n4659), .Z(n4657) );
  HS65_LS_AOI12X2 U16876 ( .A(n528), .B(n6249), .C(n6250), .Z(n6248) );
  HS65_LS_AOI12X2 U16877 ( .A(n6251), .B(n6232), .C(n6252), .Z(n6250) );
  HS65_LS_AOI12X2 U16878 ( .A(n3214), .B(n3215), .C(n2841), .Z(n3210) );
  HS65_LS_AOI12X2 U16879 ( .A(n3173), .B(n3174), .C(n2886), .Z(n3169) );
  HS65_LS_AOI12X2 U16880 ( .A(n347), .B(n8043), .C(n8044), .Z(n8042) );
  HS65_LS_AOI12X2 U16881 ( .A(n8045), .B(n8046), .C(n7952), .Z(n8044) );
  HS65_LS_AOI12X2 U16882 ( .A(n226), .B(n2963), .C(n2964), .Z(n2962) );
  HS65_LS_AOI12X2 U16883 ( .A(n2965), .B(n2945), .C(n2966), .Z(n2964) );
  HS65_LS_AOI12X2 U16884 ( .A(n2971), .B(n2972), .C(n2973), .Z(n2967) );
  HS65_LS_AOI12X2 U16885 ( .A(n3065), .B(n3066), .C(n3067), .Z(n3059) );
  HS65_LS_AOI12X2 U16886 ( .A(n7871), .B(n8009), .C(n7760), .Z(n8005) );
  HS65_LS_AOI12X2 U16887 ( .A(n7954), .B(n8051), .C(n7777), .Z(n8047) );
  HS65_LS_AOI12X2 U16888 ( .A(n7963), .B(n8332), .C(n7961), .Z(n8328) );
  HS65_LS_AOI12X2 U16889 ( .A(n7861), .B(n8136), .C(n7859), .Z(n8132) );
  HS65_LS_AOI12X2 U16890 ( .A(n2877), .B(n3133), .C(n2875), .Z(n3129) );
  HS65_LS_AOI12X2 U16891 ( .A(n177), .B(n3292), .C(n4089), .Z(n4088) );
  HS65_LS_AOI12X2 U16892 ( .A(n3067), .B(n3281), .C(n3264), .Z(n4089) );
  HS65_LS_BFX2 U16893 ( .A(n9146), .Z(n9144) );
  HS65_LS_BFX2 U16894 ( .A(n9146), .Z(n9143) );
  HS65_LS_IVX2 U16897 ( .A(n975), .Z(\u0/r0/rcnt [1]) );
  HS65_LS_BFX4 U16898 ( .A(n9148), .Z(n9147) );
  HS65_LS_IVX2 U16899 ( .A(n976), .Z(\u0/r0/rcnt [0]) );
  HS65_LS_BFX2 U16900 ( .A(n9146), .Z(n9145) );
  HS65_LS_NOR2X2 U16901 ( .A(n161), .B(n162), .Z(n4147) );
  HS65_LS_NOR2X2 U16902 ( .A(n893), .B(n892), .Z(n1478) );
  HS65_LS_NOR2X2 U16903 ( .A(n811), .B(n810), .Z(n2230) );
  HS65_LS_NOR2X2 U16904 ( .A(n934), .B(n933), .Z(n2606) );
  HS65_LS_NOR2X2 U16905 ( .A(n852), .B(n851), .Z(n1854) );
  HS65_LS_NOR2X2 U16906 ( .A(n642), .B(n651), .Z(n4281) );
  HS65_LS_NOR2X2 U16907 ( .A(n418), .B(n427), .Z(n4340) );
  HS65_LS_NOR2X2 U16908 ( .A(n333), .B(n338), .Z(n8935) );
  HS65_LS_NAND2X2 U16909 ( .A(n2595), .B(n2615), .Z(n2336) );
  HS65_LS_NAND2X2 U16910 ( .A(n1843), .B(n1863), .Z(n1584) );
  HS65_LS_NAND2X2 U16911 ( .A(n4148), .B(n4160), .Z(n3063) );
  HS65_LS_NAND2X2 U16912 ( .A(n4227), .B(n4211), .Z(n3470) );
  HS65_LS_NAND2X2 U16913 ( .A(n1467), .B(n1487), .Z(n1208) );
  HS65_LS_NAND2X2 U16914 ( .A(n4161), .B(n4148), .Z(n3045) );
  HS65_LS_NAND2X2 U16915 ( .A(n4226), .B(n4225), .Z(n3074) );
  HS65_LS_NAND2X2 U16916 ( .A(n4335), .B(n4341), .Z(n2856) );
  HS65_LS_NAND2X2 U16917 ( .A(n9029), .B(n9030), .Z(n8160) );
  HS65_LS_NAND2X2 U16918 ( .A(n9087), .B(n9088), .Z(n8192) );
  HS65_LS_NAND2X2 U16919 ( .A(n8921), .B(n8934), .Z(n8070) );
  HS65_LS_NAND2X2 U16920 ( .A(n8927), .B(n8934), .Z(n8361) );
  HS65_LS_NAND2X2 U16921 ( .A(n5748), .B(n5758), .Z(n4562) );
  HS65_LS_NAND2X2 U16922 ( .A(n7340), .B(n7350), .Z(n6155) );
  HS65_LS_NAND2X2 U16923 ( .A(n2219), .B(n2239), .Z(n1960) );
  HS65_LS_NAND2X2 U16924 ( .A(n4275), .B(n4293), .Z(n3353) );
  HS65_LS_NAND2X2 U16925 ( .A(n9057), .B(n9061), .Z(n7646) );
  HS65_LS_NAND2X2 U16926 ( .A(n9115), .B(n9119), .Z(n7674) );
  HS65_LS_NAND2X2 U16927 ( .A(n4158), .B(n4156), .Z(n3280) );
  HS65_LS_NAND2X2 U16928 ( .A(n5756), .B(n5737), .Z(n5516) );
  HS65_LS_NAND2X2 U16929 ( .A(n7348), .B(n7329), .Z(n7108) );
  HS65_LS_NAND2X2 U16930 ( .A(n5941), .B(n5940), .Z(n4509) );
  HS65_LS_NAND2X2 U16931 ( .A(n5882), .B(n5881), .Z(n4463) );
  HS65_LS_NAND2X2 U16932 ( .A(n7533), .B(n7532), .Z(n6102) );
  HS65_LS_NAND2X2 U16933 ( .A(n5815), .B(n5823), .Z(n4862) );
  HS65_LS_NAND2X2 U16934 ( .A(n7407), .B(n7415), .Z(n6455) );
  HS65_LS_NAND2X2 U16935 ( .A(n7474), .B(n7473), .Z(n6056) );
  HS65_LS_NAND2X2 U16936 ( .A(n2614), .B(n2613), .Z(n2528) );
  HS65_LS_NAND2X2 U16937 ( .A(n1862), .B(n1861), .Z(n1776) );
  HS65_LS_NAND2X2 U16938 ( .A(n1486), .B(n1485), .Z(n1400) );
  HS65_LS_NAND2X2 U16939 ( .A(n2238), .B(n2237), .Z(n2152) );
  HS65_LS_NAND2X2 U16940 ( .A(n9055), .B(n9037), .Z(n7639) );
  HS65_LS_NAND2X2 U16941 ( .A(n9113), .B(n9095), .Z(n7667) );
  HS65_LS_NAND2X2 U16942 ( .A(n5754), .B(n5751), .Z(n4560) );
  HS65_LS_NAND2X2 U16943 ( .A(n7346), .B(n7343), .Z(n6153) );
  HS65_LS_NAND2X2 U16944 ( .A(n4211), .B(n4230), .Z(n2965) );
  HS65_LS_NAND2X2 U16945 ( .A(n5934), .B(n5946), .Z(n4511) );
  HS65_LS_NAND2X2 U16946 ( .A(n5875), .B(n5887), .Z(n4465) );
  HS65_LS_NAND2X2 U16947 ( .A(n7526), .B(n7538), .Z(n6104) );
  HS65_LS_NAND2X2 U16948 ( .A(n7467), .B(n7479), .Z(n6058) );
  HS65_LS_NAND2X2 U16949 ( .A(n5816), .B(n5813), .Z(n4636) );
  HS65_LS_NAND2X2 U16950 ( .A(n7408), .B(n7405), .Z(n6229) );
  HS65_LS_NAND2X2 U16951 ( .A(n4349), .B(n4348), .Z(n3983) );
  HS65_LS_NAND2X2 U16952 ( .A(n4337), .B(n4351), .Z(n3895) );
  HS65_LS_NAND2X2 U16953 ( .A(n8988), .B(n8987), .Z(n8220) );
  HS65_LS_NAND2X2 U16954 ( .A(n4161), .B(n4150), .Z(n2927) );
  HS65_LS_NAND2X2 U16955 ( .A(n9095), .B(n9096), .Z(n8182) );
  HS65_LS_NAND2X2 U16956 ( .A(n9037), .B(n9038), .Z(n8150) );
  HS65_LS_NAND2X2 U16957 ( .A(n9053), .B(n9044), .Z(n8412) );
  HS65_LS_NAND2X2 U16958 ( .A(n9111), .B(n9102), .Z(n8472) );
  HS65_LS_NAND2X2 U16959 ( .A(n8929), .B(n8918), .Z(n8045) );
  HS65_LS_NAND2X2 U16960 ( .A(n4226), .B(n4229), .Z(n3536) );
  HS65_LS_NAND2X2 U16961 ( .A(n5756), .B(n5757), .Z(n4577) );
  HS65_LS_NAND2X2 U16962 ( .A(n7348), .B(n7349), .Z(n6170) );
  HS65_LS_NAND2X2 U16963 ( .A(n5939), .B(n5920), .Z(n5639) );
  HS65_LS_NAND2X2 U16964 ( .A(n5880), .B(n5861), .Z(n5612) );
  HS65_LS_NAND2X2 U16965 ( .A(n7531), .B(n7512), .Z(n7231) );
  HS65_LS_NAND2X2 U16966 ( .A(n7472), .B(n7453), .Z(n7204) );
  HS65_LS_NAND2X2 U16967 ( .A(n5818), .B(n5814), .Z(n5588) );
  HS65_LS_NAND2X2 U16968 ( .A(n7410), .B(n7406), .Z(n7180) );
  HS65_LS_NAND2X2 U16969 ( .A(n4158), .B(n4168), .Z(n3264) );
  HS65_LS_NAND2X2 U16970 ( .A(n9037), .B(n9051), .Z(n7818) );
  HS65_LS_NAND2X2 U16971 ( .A(n9095), .B(n9109), .Z(n7917) );
  HS65_LS_NAND2X2 U16972 ( .A(n2592), .B(n2595), .Z(n2504) );
  HS65_LS_NAND2X2 U16973 ( .A(n1464), .B(n1467), .Z(n1376) );
  HS65_LS_NAND2X2 U16974 ( .A(n2216), .B(n2219), .Z(n2128) );
  HS65_LS_NAND2X2 U16975 ( .A(n1840), .B(n1843), .Z(n1752) );
  HS65_LS_NOR2X2 U16976 ( .A(n405), .B(n406), .Z(n8997) );
  HS65_LS_NAND2X2 U16977 ( .A(n4150), .B(n4160), .Z(n2923) );
  HS65_LS_NAND2X2 U16978 ( .A(n8994), .B(n9001), .Z(n8095) );
  HS65_LS_NAND2X2 U16979 ( .A(n4155), .B(n4156), .Z(n3043) );
  HS65_LS_NAND2X2 U16980 ( .A(n7467), .B(n7477), .Z(n6353) );
  HS65_LS_NAND2X2 U16981 ( .A(n5934), .B(n5944), .Z(n4799) );
  HS65_LS_NAND2X2 U16982 ( .A(n7526), .B(n7536), .Z(n6392) );
  HS65_LS_NAND2X2 U16983 ( .A(n5875), .B(n5885), .Z(n4760) );
  HS65_LS_NAND2X2 U16984 ( .A(n5816), .B(n5817), .Z(n4653) );
  HS65_LS_NAND2X2 U16985 ( .A(n7408), .B(n7409), .Z(n6246) );
  HS65_LS_NAND2X2 U16986 ( .A(n7352), .B(n7353), .Z(n7109) );
  HS65_LS_NAND2X2 U16987 ( .A(n5760), .B(n5761), .Z(n5517) );
  HS65_LS_NAND2X2 U16988 ( .A(n5754), .B(n5755), .Z(n4576) );
  HS65_LS_NAND2X2 U16989 ( .A(n7346), .B(n7347), .Z(n6169) );
  HS65_LS_NAND2X2 U16990 ( .A(n4227), .B(n4222), .Z(n2943) );
  HS65_LS_NAND2X2 U16991 ( .A(n7453), .B(n7454), .Z(n6488) );
  HS65_LS_NAND2X2 U16992 ( .A(n5861), .B(n5862), .Z(n4895) );
  HS65_LS_NAND2X2 U16993 ( .A(n5920), .B(n5921), .Z(n5009) );
  HS65_LS_NAND2X2 U16994 ( .A(n7512), .B(n7513), .Z(n6602) );
  HS65_LS_NAND2X2 U16995 ( .A(n7344), .B(n7330), .Z(n6270) );
  HS65_LS_NAND2X2 U16996 ( .A(n5752), .B(n5738), .Z(n4677) );
  HS65_LS_NAND2X2 U16997 ( .A(n5814), .B(n5800), .Z(n4881) );
  HS65_LS_NAND2X2 U16998 ( .A(n7406), .B(n7392), .Z(n6474) );
  HS65_LS_NAND2X2 U16999 ( .A(n9001), .B(n9002), .Z(n8009) );
  HS65_LS_NAND2X2 U17000 ( .A(n4161), .B(n4162), .Z(n3625) );
  HS65_LS_NOR2X2 U17001 ( .A(n871), .B(n870), .Z(n1465) );
  HS65_LS_NOR2X2 U17002 ( .A(n789), .B(n788), .Z(n2217) );
  HS65_LS_NOR2X2 U17003 ( .A(n830), .B(n829), .Z(n1841) );
  HS65_LS_NOR2X2 U17004 ( .A(n912), .B(n911), .Z(n2593) );
  HS65_LS_NAND2X2 U17005 ( .A(n2596), .B(n2603), .Z(n2282) );
  HS65_LS_NAND2X2 U17006 ( .A(n1844), .B(n1851), .Z(n1530) );
  HS65_LS_NAND2X2 U17007 ( .A(n4279), .B(n4280), .Z(n2895) );
  HS65_LS_NAND2X2 U17008 ( .A(n4294), .B(n4274), .Z(n3726) );
  HS65_LS_NAND2X2 U17009 ( .A(n9054), .B(n9061), .Z(n7832) );
  HS65_LS_NAND2X2 U17010 ( .A(n9112), .B(n9119), .Z(n7931) );
  HS65_LS_NAND2X2 U17011 ( .A(n1468), .B(n1475), .Z(n1154) );
  HS65_LS_NAND2X2 U17012 ( .A(n2220), .B(n2227), .Z(n1906) );
  HS65_LS_NAND2X2 U17013 ( .A(n9113), .B(n9114), .Z(n7663) );
  HS65_LS_NAND2X2 U17014 ( .A(n9055), .B(n9056), .Z(n7635) );
  HS65_LS_NAND2X2 U17015 ( .A(n5755), .B(n5762), .Z(n5492) );
  HS65_LS_NAND2X2 U17016 ( .A(n7347), .B(n7354), .Z(n7084) );
  HS65_LS_NAND2X2 U17017 ( .A(n1866), .B(n1852), .Z(n1686) );
  HS65_LS_NAND2X2 U17018 ( .A(n2618), .B(n2604), .Z(n2438) );
  HS65_LS_NAND2X2 U17019 ( .A(n5944), .B(n5945), .Z(n4517) );
  HS65_LS_NAND2X2 U17020 ( .A(n5885), .B(n5886), .Z(n4471) );
  HS65_LS_NAND2X2 U17021 ( .A(n7536), .B(n7537), .Z(n6110) );
  HS65_LS_NAND2X2 U17022 ( .A(n5817), .B(n5824), .Z(n5508) );
  HS65_LS_NAND2X2 U17023 ( .A(n7409), .B(n7416), .Z(n7100) );
  HS65_LS_NAND2X2 U17024 ( .A(n7477), .B(n7478), .Z(n6064) );
  HS65_LS_NAND2X2 U17025 ( .A(n4227), .B(n4213), .Z(n2873) );
  HS65_LS_NAND2X2 U17026 ( .A(n4169), .B(n4161), .Z(n3599) );
  HS65_LS_NAND2X2 U17027 ( .A(n1490), .B(n1476), .Z(n1310) );
  HS65_LS_NAND2X2 U17028 ( .A(n4276), .B(n4282), .Z(n2901) );
  HS65_LS_NAND2X2 U17029 ( .A(n4277), .B(n4290), .Z(n3147) );
  HS65_LS_NAND2X2 U17030 ( .A(n8981), .B(n9002), .Z(n8031) );
  HS65_LS_NAND2X2 U17031 ( .A(n5753), .B(n5737), .Z(n5039) );
  HS65_LS_NAND2X2 U17032 ( .A(n7345), .B(n7329), .Z(n6632) );
  HS65_LS_NAND2X2 U17033 ( .A(n5941), .B(n5931), .Z(n5393) );
  HS65_LS_NAND2X2 U17034 ( .A(n5882), .B(n5872), .Z(n5278) );
  HS65_LS_NAND2X2 U17035 ( .A(n5815), .B(n5799), .Z(n5161) );
  HS65_LS_NAND2X2 U17036 ( .A(n7533), .B(n7523), .Z(n6985) );
  HS65_LS_NAND2X2 U17037 ( .A(n7407), .B(n7391), .Z(n6753) );
  HS65_LS_NAND2X2 U17038 ( .A(n7474), .B(n7464), .Z(n6870) );
  HS65_LS_NAND2X2 U17039 ( .A(n4222), .B(n4230), .Z(n2960) );
  HS65_LS_NAND2X2 U17040 ( .A(n2242), .B(n2228), .Z(n2062) );
  HS65_LS_NAND2X2 U17041 ( .A(n8988), .B(n8978), .Z(n8004) );
  HS65_LS_NAND2X2 U17042 ( .A(n7456), .B(n7466), .Z(n6339) );
  HS65_LS_NAND2X2 U17043 ( .A(n5923), .B(n5933), .Z(n4785) );
  HS65_LS_NAND2X2 U17044 ( .A(n7515), .B(n7525), .Z(n6378) );
  HS65_LS_NAND2X2 U17045 ( .A(n5864), .B(n5874), .Z(n4746) );
  HS65_LS_NAND2X2 U17046 ( .A(n5810), .B(n5820), .Z(n4639) );
  HS65_LS_NAND2X2 U17047 ( .A(n7402), .B(n7412), .Z(n6232) );
  HS65_LS_NAND2X2 U17048 ( .A(n5760), .B(n5757), .Z(n4669) );
  HS65_LS_NAND2X2 U17049 ( .A(n7352), .B(n7349), .Z(n6262) );
  HS65_LS_NAND2X2 U17050 ( .A(n7454), .B(n7473), .Z(n6065) );
  HS65_LS_NAND2X2 U17051 ( .A(n7513), .B(n7532), .Z(n6111) );
  HS65_LS_NAND2X2 U17052 ( .A(n5862), .B(n5881), .Z(n4472) );
  HS65_LS_NAND2X2 U17053 ( .A(n5921), .B(n5940), .Z(n4518) );
  HS65_LS_NAND2X2 U17054 ( .A(n5800), .B(n5823), .Z(n4533) );
  HS65_LS_NAND2X2 U17055 ( .A(n7392), .B(n7415), .Z(n6126) );
  HS65_LS_NAND2X2 U17056 ( .A(n7472), .B(n7464), .Z(n7137) );
  HS65_LS_NAND2X2 U17057 ( .A(n5939), .B(n5931), .Z(n5566) );
  HS65_LS_NAND2X2 U17058 ( .A(n7531), .B(n7523), .Z(n7158) );
  HS65_LS_NAND2X2 U17059 ( .A(n5880), .B(n5872), .Z(n5545) );
  HS65_LS_NAND2X2 U17060 ( .A(n5818), .B(n5799), .Z(n5581) );
  HS65_LS_NAND2X2 U17061 ( .A(n7410), .B(n7391), .Z(n7173) );
  HS65_LS_NAND2X2 U17062 ( .A(n4338), .B(n4337), .Z(n3003) );
  HS65_LS_NAND2X2 U17063 ( .A(n4226), .B(n4219), .Z(n3102) );
  HS65_LS_NAND2X2 U17064 ( .A(n4157), .B(n4165), .Z(n4002) );
  HS65_LS_NOR2X2 U17065 ( .A(n339), .B(n340), .Z(n8928) );
  HS65_LS_NOR2X2 U17066 ( .A(n382), .B(n383), .Z(n8998) );
  HS65_LS_NOR2X2 U17067 ( .A(n429), .B(n428), .Z(n4339) );
  HS65_LS_NOR2X2 U17068 ( .A(n603), .B(n602), .Z(n9053) );
  HS65_LS_NOR2X2 U17069 ( .A(n116), .B(n115), .Z(n9111) );
  HS65_LS_NOR2X2 U17070 ( .A(n206), .B(n207), .Z(n4212) );
  HS65_LS_NOR2X2 U17071 ( .A(n117), .B(n118), .Z(n9088) );
  HS65_LS_NOR2X2 U17072 ( .A(n604), .B(n605), .Z(n9030) );
  HS65_LS_NOR2X2 U17073 ( .A(n360), .B(n361), .Z(n8942) );
  HS65_LS_NOR2X2 U17074 ( .A(n449), .B(n450), .Z(n4341) );
  HS65_LS_NOR2X2 U17075 ( .A(n229), .B(n230), .Z(n4225) );
  HS65_LS_NAND2X2 U17076 ( .A(n4333), .B(n4348), .Z(n3215) );
  HS65_LS_NAND2X2 U17077 ( .A(n4290), .B(n4287), .Z(n3167) );
  HS65_LS_NAND2X2 U17078 ( .A(n1468), .B(n1469), .Z(n1130) );
  HS65_LS_NAND2X2 U17079 ( .A(n2220), .B(n2221), .Z(n1882) );
  HS65_LS_NAND2X2 U17080 ( .A(n2596), .B(n2597), .Z(n2258) );
  HS65_LS_NAND2X2 U17081 ( .A(n1844), .B(n1845), .Z(n1506) );
  HS65_LS_NAND2X2 U17082 ( .A(n1850), .B(n1865), .Z(n1529) );
  HS65_LS_NAND2X2 U17083 ( .A(n2602), .B(n2617), .Z(n2281) );
  HS65_LS_NAND2X2 U17084 ( .A(n4157), .B(n4158), .Z(n3058) );
  HS65_LS_NAND2X2 U17085 ( .A(n7347), .B(n7342), .Z(n7118) );
  HS65_LS_NAND2X2 U17086 ( .A(n5755), .B(n5750), .Z(n5526) );
  HS65_LS_NAND2X2 U17087 ( .A(n7472), .B(n7476), .Z(n6354) );
  HS65_LS_NAND2X2 U17088 ( .A(n5939), .B(n5943), .Z(n4800) );
  HS65_LS_NAND2X2 U17089 ( .A(n7531), .B(n7535), .Z(n6393) );
  HS65_LS_NAND2X2 U17090 ( .A(n5880), .B(n5884), .Z(n4761) );
  HS65_LS_NAND2X2 U17091 ( .A(n5818), .B(n5819), .Z(n4654) );
  HS65_LS_NAND2X2 U17092 ( .A(n7410), .B(n7411), .Z(n6247) );
  HS65_LS_NAND2X2 U17093 ( .A(n4168), .B(n4165), .Z(n3064) );
  HS65_LS_NAND2X2 U17094 ( .A(n9000), .B(n8978), .Z(n8003) );
  HS65_LS_NAND2X2 U17095 ( .A(n9050), .B(n9059), .Z(n8436) );
  HS65_LS_NAND2X2 U17096 ( .A(n9108), .B(n9117), .Z(n8447) );
  HS65_LS_NAND2X2 U17097 ( .A(n1474), .B(n1489), .Z(n1153) );
  HS65_LS_NAND2X2 U17098 ( .A(n2226), .B(n2241), .Z(n1905) );
  HS65_LS_NAND2X2 U17099 ( .A(n5756), .B(n5752), .Z(n5523) );
  HS65_LS_NAND2X2 U17100 ( .A(n7348), .B(n7344), .Z(n7115) );
  HS65_LS_NAND2X2 U17101 ( .A(n9109), .B(n9114), .Z(n7893) );
  HS65_LS_NAND2X2 U17102 ( .A(n9051), .B(n9056), .Z(n7793) );
  HS65_LS_NAND2X2 U17103 ( .A(n4231), .B(n4224), .Z(n2961) );
  HS65_LS_NAND2X2 U17104 ( .A(n4155), .B(n4168), .Z(n3236) );
  HS65_LS_NAND2X2 U17105 ( .A(n4221), .B(n4228), .Z(n3454) );
  HS65_LS_NAND2X2 U17106 ( .A(n4336), .B(n4352), .Z(n3002) );
  HS65_LS_NAND2X2 U17107 ( .A(n4277), .B(n4288), .Z(n2984) );
  HS65_LS_NAND2X2 U17108 ( .A(n8926), .B(n8927), .Z(n8542) );
  HS65_LS_NAND2X2 U17109 ( .A(n2602), .B(n2612), .Z(n2300) );
  HS65_LS_NAND2X2 U17110 ( .A(n1850), .B(n1860), .Z(n1548) );
  HS65_LS_NAND2X2 U17111 ( .A(n4160), .B(n4162), .Z(n3042) );
  HS65_LS_NAND2X2 U17112 ( .A(n1474), .B(n1484), .Z(n1172) );
  HS65_LS_NAND2X2 U17113 ( .A(n2226), .B(n2236), .Z(n1924) );
  HS65_LS_NAND2X2 U17114 ( .A(n5756), .B(n5761), .Z(n4695) );
  HS65_LS_NAND2X2 U17115 ( .A(n7348), .B(n7353), .Z(n6288) );
  HS65_LS_NAND2X2 U17116 ( .A(n8994), .B(n8997), .Z(n8080) );
  HS65_LS_NAND2X2 U17117 ( .A(n4336), .B(n4347), .Z(n3188) );
  HS65_LS_NAND2X2 U17118 ( .A(n5933), .B(n5945), .Z(n4620) );
  HS65_LS_NAND2X2 U17119 ( .A(n5874), .B(n5886), .Z(n4595) );
  HS65_LS_NAND2X2 U17120 ( .A(n7525), .B(n7537), .Z(n6213) );
  HS65_LS_NAND2X2 U17121 ( .A(n5820), .B(n5824), .Z(n5148) );
  HS65_LS_NAND2X2 U17122 ( .A(n5758), .B(n5762), .Z(n5026) );
  HS65_LS_NAND2X2 U17123 ( .A(n7466), .B(n7478), .Z(n6188) );
  HS65_LS_NAND2X2 U17124 ( .A(n7350), .B(n7354), .Z(n6619) );
  HS65_LS_NAND2X2 U17125 ( .A(n7412), .B(n7416), .Z(n6740) );
  HS65_LS_NAND2X2 U17126 ( .A(n4167), .B(n4163), .Z(n3290) );
  HS65_LS_NAND2X2 U17127 ( .A(n4167), .B(n4168), .Z(n3585) );
  HS65_LS_NAND2X2 U17128 ( .A(n4279), .B(n4278), .Z(n2985) );
  HS65_LS_NAND2X2 U17129 ( .A(n8926), .B(n8942), .Z(n8335) );
  HS65_LS_NAND2X2 U17130 ( .A(n4349), .B(n4334), .Z(n3985) );
  HS65_LS_NAND2X2 U17131 ( .A(n8920), .B(n8940), .Z(n8041) );
  HS65_LS_NAND2X2 U17132 ( .A(n4280), .B(n4287), .Z(n3162) );
  HS65_LS_NAND2X2 U17133 ( .A(n4219), .B(n4223), .Z(n3484) );
  HS65_LS_NAND2X2 U17134 ( .A(n4353), .B(n4333), .Z(n3843) );
  HS65_LS_NAND2X2 U17135 ( .A(n8939), .B(n8918), .Z(n8046) );
  HS65_LS_NAND2X2 U17136 ( .A(n7463), .B(n7476), .Z(n6481) );
  HS65_LS_NAND2X2 U17137 ( .A(n7522), .B(n7535), .Z(n6595) );
  HS65_LS_NAND2X2 U17138 ( .A(n5871), .B(n5884), .Z(n4888) );
  HS65_LS_NAND2X2 U17139 ( .A(n5930), .B(n5943), .Z(n5002) );
  HS65_LS_NAND2X2 U17140 ( .A(n5822), .B(n5819), .Z(n4874) );
  HS65_LS_NAND2X2 U17141 ( .A(n7414), .B(n7411), .Z(n6467) );
  HS65_LS_NAND2X2 U17142 ( .A(n8999), .B(n9000), .Z(n7998) );
  HS65_LS_NAND2X2 U17143 ( .A(n4292), .B(n4291), .Z(n3962) );
  HS65_LS_NAND2X2 U17144 ( .A(n4335), .B(n4353), .Z(n2847) );
  HS65_LS_NAND2X2 U17145 ( .A(n4276), .B(n4294), .Z(n2892) );
  HS65_LS_NAND2X2 U17146 ( .A(n4221), .B(n4211), .Z(n2945) );
  HS65_LS_NAND2X2 U17147 ( .A(n2242), .B(n2238), .Z(n1953) );
  HS65_LS_NAND2X2 U17148 ( .A(n1866), .B(n1862), .Z(n1577) );
  HS65_LS_NAND2X2 U17149 ( .A(n2618), .B(n2614), .Z(n2329) );
  HS65_LS_NAND2X2 U17150 ( .A(n1490), .B(n1486), .Z(n1201) );
  HS65_LS_NAND2X2 U17151 ( .A(n4292), .B(n4275), .Z(n3964) );
  HS65_LS_NAND2X2 U17152 ( .A(n4220), .B(n4229), .Z(n3942) );
  HS65_LS_NOR2X2 U17153 ( .A(n890), .B(n891), .Z(n1469) );
  HS65_LS_NOR2X2 U17154 ( .A(n808), .B(n809), .Z(n2221) );
  HS65_LS_NOR2X2 U17155 ( .A(n931), .B(n932), .Z(n2597) );
  HS65_LS_NOR2X2 U17156 ( .A(n849), .B(n850), .Z(n1845) );
  HS65_LS_NAND2X2 U17157 ( .A(n4293), .B(n4291), .Z(n3163) );
  HS65_LS_NAND2X2 U17158 ( .A(n9057), .B(n9029), .Z(n8164) );
  HS65_LS_NAND2X2 U17159 ( .A(n9115), .B(n9087), .Z(n8196) );
  HS65_LS_NAND2X2 U17160 ( .A(n7477), .B(n7465), .Z(n7210) );
  HS65_LS_NAND2X2 U17161 ( .A(n5944), .B(n5932), .Z(n5645) );
  HS65_LS_NAND2X2 U17162 ( .A(n7536), .B(n7524), .Z(n7237) );
  HS65_LS_NAND2X2 U17163 ( .A(n5885), .B(n5873), .Z(n5618) );
  HS65_LS_NAND2X2 U17164 ( .A(n5817), .B(n5812), .Z(n5591) );
  HS65_LS_NAND2X2 U17165 ( .A(n7409), .B(n7404), .Z(n7183) );
  HS65_LS_NAND2X2 U17166 ( .A(n4220), .B(n4224), .Z(n3940) );
  HS65_LS_NAND2X2 U17167 ( .A(n2615), .B(n2613), .Z(n2324) );
  HS65_LS_NAND2X2 U17168 ( .A(n1863), .B(n1861), .Z(n1572) );
  HS65_LS_NAND2X2 U17169 ( .A(n7330), .B(n7353), .Z(n6086) );
  HS65_LS_NAND2X2 U17170 ( .A(n5738), .B(n5761), .Z(n4493) );
  HS65_LS_NAND2X2 U17171 ( .A(n9050), .B(n9038), .Z(n7644) );
  HS65_LS_NAND2X2 U17172 ( .A(n9108), .B(n9096), .Z(n7672) );
  HS65_LS_NAND2X2 U17173 ( .A(n5752), .B(n5753), .Z(n4582) );
  HS65_LS_NAND2X2 U17174 ( .A(n7344), .B(n7345), .Z(n6175) );
  HS65_LS_NAND2X2 U17175 ( .A(n1486), .B(n1467), .Z(n1404) );
  HS65_LS_NAND2X2 U17176 ( .A(n2238), .B(n2219), .Z(n2156) );
  HS65_LS_NAND2X2 U17177 ( .A(n1862), .B(n1843), .Z(n1780) );
  HS65_LS_NAND2X2 U17178 ( .A(n2614), .B(n2595), .Z(n2532) );
  HS65_LS_NAND2X2 U17179 ( .A(n8980), .B(n9001), .Z(n7999) );
  HS65_LS_NAND2X2 U17180 ( .A(n1487), .B(n1485), .Z(n1196) );
  HS65_LS_NAND2X2 U17181 ( .A(n2239), .B(n2237), .Z(n1948) );
  HS65_LS_NAND2X2 U17182 ( .A(n8996), .B(n8981), .Z(n7869) );
  HS65_LS_NAND2X2 U17183 ( .A(n4350), .B(n4348), .Z(n3204) );
  HS65_LS_NAND2X2 U17184 ( .A(n2597), .B(n2616), .Z(n2323) );
  HS65_LS_NAND2X2 U17185 ( .A(n1845), .B(n1864), .Z(n1571) );
  HS65_LS_NAND2X2 U17186 ( .A(n1469), .B(n1488), .Z(n1195) );
  HS65_LS_NAND2X2 U17187 ( .A(n2221), .B(n2240), .Z(n1947) );
  HS65_LS_NAND2X2 U17188 ( .A(n9052), .B(n9051), .Z(n7633) );
  HS65_LS_NAND2X2 U17189 ( .A(n9110), .B(n9109), .Z(n7661) );
  HS65_LS_NAND2X2 U17190 ( .A(n1852), .B(n1861), .Z(n1777) );
  HS65_LS_NAND2X2 U17191 ( .A(n2604), .B(n2613), .Z(n2529) );
  HS65_LS_NAND2X2 U17192 ( .A(n4157), .B(n4167), .Z(n4103) );
  HS65_LS_NOR2X2 U17193 ( .A(n672), .B(n673), .Z(n4276) );
  HS65_LS_NAND2X2 U17194 ( .A(n2228), .B(n2237), .Z(n2153) );
  HS65_LS_NAND2X2 U17195 ( .A(n1476), .B(n1485), .Z(n1401) );
  HS65_LS_NOR2X2 U17196 ( .A(n384), .B(n385), .Z(n8999) );
  HS65_LS_NOR2X2 U17197 ( .A(n653), .B(n652), .Z(n4280) );
  HS65_LS_NAND2X2 U17198 ( .A(n4223), .B(n4224), .Z(n2972) );
  HS65_LS_NOR2X2 U17199 ( .A(n134), .B(n139), .Z(n9114) );
  HS65_LS_NOR2X2 U17200 ( .A(n621), .B(n626), .Z(n9056) );
  HS65_LS_NOR2X2 U17201 ( .A(n490), .B(n491), .Z(n5940) );
  HS65_LS_NOR2X2 U17202 ( .A(n271), .B(n272), .Z(n5881) );
  HS65_LS_NOR2X2 U17203 ( .A(n313), .B(n314), .Z(n7532) );
  HS65_LS_NOR2X2 U17204 ( .A(n92), .B(n93), .Z(n7473) );
  HS65_LS_NOR2X2 U17205 ( .A(n708), .B(n713), .Z(n5823) );
  HS65_LS_NOR2X2 U17206 ( .A(n526), .B(n531), .Z(n7415) );
  HS65_LS_NAND2X2 U17207 ( .A(n8996), .B(n8995), .Z(n8671) );
  HS65_LS_NAND2X2 U17208 ( .A(n8928), .B(n8929), .Z(n8040) );
  HS65_LS_NAND2X2 U17209 ( .A(n4339), .B(n4351), .Z(n3203) );
  HS65_LS_NAND2X2 U17210 ( .A(n1464), .B(n1490), .Z(n1127) );
  HS65_LS_NAND2X2 U17211 ( .A(n1840), .B(n1866), .Z(n1503) );
  HS65_LS_NAND2X2 U17212 ( .A(n2592), .B(n2618), .Z(n2255) );
  HS65_LS_NAND2X2 U17213 ( .A(n2216), .B(n2242), .Z(n1879) );
  HS65_LS_NAND2X2 U17214 ( .A(n8941), .B(n8921), .Z(n7952) );
  HS65_LS_NAND2X2 U17215 ( .A(n4219), .B(n4220), .Z(n2966) );
  HS65_LS_NAND2X2 U17216 ( .A(n4353), .B(n4349), .Z(n3209) );
  HS65_LS_NAND2X2 U17217 ( .A(n4164), .B(n4162), .Z(n3052) );
  HS65_LS_NAND2X2 U17218 ( .A(n7477), .B(n7456), .Z(n6358) );
  HS65_LS_NAND2X2 U17219 ( .A(n5944), .B(n5923), .Z(n4804) );
  HS65_LS_NAND2X2 U17220 ( .A(n7536), .B(n7515), .Z(n6397) );
  HS65_LS_NAND2X2 U17221 ( .A(n5885), .B(n5864), .Z(n4765) );
  HS65_LS_NAND2X2 U17222 ( .A(n5817), .B(n5810), .Z(n4658) );
  HS65_LS_NAND2X2 U17223 ( .A(n7409), .B(n7402), .Z(n6251) );
  HS65_LS_NAND2X2 U17224 ( .A(n8941), .B(n8927), .Z(n8881) );
  HS65_LS_NAND2X2 U17225 ( .A(n5920), .B(n5941), .Z(n4805) );
  HS65_LS_NAND2X2 U17226 ( .A(n7512), .B(n7533), .Z(n6398) );
  HS65_LS_NAND2X2 U17227 ( .A(n7453), .B(n7474), .Z(n6359) );
  HS65_LS_NAND2X2 U17228 ( .A(n5861), .B(n5882), .Z(n4766) );
  HS65_LS_NAND2X2 U17229 ( .A(n7406), .B(n7407), .Z(n6252) );
  HS65_LS_NAND2X2 U17230 ( .A(n5814), .B(n5815), .Z(n4659) );
  HS65_LS_NOR2X2 U17231 ( .A(n873), .B(n872), .Z(n1464) );
  HS65_LS_NOR2X2 U17232 ( .A(n914), .B(n913), .Z(n2592) );
  HS65_LS_NOR2X2 U17233 ( .A(n832), .B(n831), .Z(n1840) );
  HS65_LS_NOR2X2 U17234 ( .A(n791), .B(n790), .Z(n2216) );
  HS65_LS_NAND2X2 U17235 ( .A(n9055), .B(n9050), .Z(n7978) );
  HS65_LS_NAND2X2 U17236 ( .A(n9113), .B(n9108), .Z(n7991) );
  HS65_LS_NAND2X2 U17237 ( .A(n7352), .B(n7344), .Z(n6087) );
  HS65_LS_NAND2X2 U17238 ( .A(n5760), .B(n5752), .Z(n4494) );
  HS65_LS_NAND2X2 U17239 ( .A(n4225), .B(n4231), .Z(n2971) );
  HS65_LS_NAND2X2 U17240 ( .A(n5930), .B(n5920), .Z(n4618) );
  HS65_LS_NAND2X2 U17241 ( .A(n7522), .B(n7512), .Z(n6211) );
  HS65_LS_NAND2X2 U17242 ( .A(n7463), .B(n7453), .Z(n6186) );
  HS65_LS_NAND2X2 U17243 ( .A(n5871), .B(n5861), .Z(n4593) );
  HS65_LS_NAND2X2 U17244 ( .A(n5822), .B(n5814), .Z(n4534) );
  HS65_LS_NAND2X2 U17245 ( .A(n7414), .B(n7406), .Z(n6127) );
  HS65_LS_NAND2X2 U17246 ( .A(n4337), .B(n4340), .Z(n3004) );
  HS65_LS_NAND2X2 U17247 ( .A(n8998), .B(n8989), .Z(n7858) );
  HS65_LS_NAND2X2 U17248 ( .A(n8935), .B(n8936), .Z(n7960) );
  HS65_LS_NAND2X2 U17249 ( .A(n8942), .B(n8920), .Z(n7954) );
  HS65_LS_NAND2X2 U17250 ( .A(n4338), .B(n4352), .Z(n2841) );
  HS65_LS_NAND2X2 U17251 ( .A(n4279), .B(n4288), .Z(n2886) );
  HS65_LS_NAND2X2 U17252 ( .A(n4278), .B(n4281), .Z(n2986) );
  HS65_LS_NAND2X2 U17253 ( .A(n4294), .B(n4292), .Z(n3168) );
  HS65_LS_NAND2X2 U17254 ( .A(n4341), .B(n4350), .Z(n3214) );
  HS65_LS_NAND2X2 U17255 ( .A(n5755), .B(n5748), .Z(n4581) );
  HS65_LS_NAND2X2 U17256 ( .A(n7347), .B(n7340), .Z(n6174) );
  HS65_LS_NAND2X2 U17257 ( .A(n4155), .B(n4163), .Z(n3065) );
  HS65_LS_NAND2X2 U17258 ( .A(n9054), .B(n9058), .Z(n7686) );
  HS65_LS_NAND2X2 U17259 ( .A(n9112), .B(n9116), .Z(n7724) );
  HS65_LS_NOR2X2 U17260 ( .A(n209), .B(n208), .Z(n4222) );
  HS65_LS_NAND2X2 U17261 ( .A(n1844), .B(n1865), .Z(n1497) );
  HS65_LS_NAND2X2 U17262 ( .A(n2596), .B(n2617), .Z(n2249) );
  HS65_LS_NAND2X2 U17263 ( .A(n2227), .B(n2230), .Z(n1907) );
  HS65_LS_NAND2X2 U17264 ( .A(n1475), .B(n1478), .Z(n1155) );
  HS65_LS_NAND2X2 U17265 ( .A(n2603), .B(n2606), .Z(n2283) );
  HS65_LS_NAND2X2 U17266 ( .A(n1851), .B(n1854), .Z(n1531) );
  HS65_LS_NOR2X2 U17267 ( .A(n44), .B(n49), .Z(n5761) );
  HS65_LS_NOR2X2 U17268 ( .A(n570), .B(n575), .Z(n7353) );
  HS65_LS_NOR2X2 U17269 ( .A(n163), .B(n164), .Z(n4162) );
  HS65_LS_NAND2X2 U17270 ( .A(n2220), .B(n2241), .Z(n1873) );
  HS65_LS_NAND2X2 U17271 ( .A(n1468), .B(n1489), .Z(n1121) );
  HS65_LS_NAND2X2 U17272 ( .A(n4213), .B(n4212), .Z(n2874) );
  HS65_LS_NAND2X2 U17273 ( .A(n8928), .B(n8917), .Z(n7955) );
  HS65_LS_NAND2X2 U17274 ( .A(n5750), .B(n5749), .Z(n4720) );
  HS65_LS_NAND2X2 U17275 ( .A(n7342), .B(n7341), .Z(n6313) );
  HS65_LS_NAND2X2 U17276 ( .A(n5932), .B(n5924), .Z(n4989) );
  HS65_LS_NAND2X2 U17277 ( .A(n7524), .B(n7516), .Z(n6582) );
  HS65_LS_NAND2X2 U17278 ( .A(n7465), .B(n7457), .Z(n6528) );
  HS65_LS_NAND2X2 U17279 ( .A(n5873), .B(n5865), .Z(n4935) );
  HS65_LS_NAND2X2 U17280 ( .A(n7404), .B(n7403), .Z(n6452) );
  HS65_LS_NAND2X2 U17281 ( .A(n5812), .B(n5811), .Z(n4859) );
  HS65_LS_NAND2X2 U17282 ( .A(n4282), .B(n4293), .Z(n3173) );
  HS65_LS_NAND2X2 U17283 ( .A(n7479), .B(n7478), .Z(n6051) );
  HS65_LS_NAND2X2 U17284 ( .A(n7405), .B(n7416), .Z(n6413) );
  HS65_LS_NAND2X2 U17285 ( .A(n5813), .B(n5824), .Z(n4820) );
  HS65_LS_NAND2X2 U17286 ( .A(n5946), .B(n5945), .Z(n4504) );
  HS65_LS_NAND2X2 U17287 ( .A(n7538), .B(n7537), .Z(n6097) );
  HS65_LS_NAND2X2 U17288 ( .A(n5887), .B(n5886), .Z(n4458) );
  HS65_LS_NAND2X2 U17289 ( .A(n8988), .B(n8989), .Z(n7861) );
  HS65_LS_NAND2X2 U17290 ( .A(n8939), .B(n8936), .Z(n7963) );
  HS65_LS_NAND2X2 U17291 ( .A(n4227), .B(n4228), .Z(n2973) );
  HS65_LS_NAND2X2 U17292 ( .A(n5751), .B(n5762), .Z(n4680) );
  HS65_LS_NAND2X2 U17293 ( .A(n7343), .B(n7354), .Z(n6273) );
  HS65_LS_NAND2X2 U17294 ( .A(n4333), .B(n4334), .Z(n2849) );
  HS65_LS_NAND2X2 U17295 ( .A(n8941), .B(n8940), .Z(n8639) );
  HS65_LS_NAND2X2 U17296 ( .A(n8935), .B(n8938), .Z(n8332) );
  HS65_LS_NAND2X2 U17297 ( .A(n4228), .B(n4212), .Z(n3133) );
  HS65_LS_NAND2X2 U17298 ( .A(n4288), .B(n4281), .Z(n3359) );
  HS65_LS_NAND2X2 U17299 ( .A(n4352), .B(n4340), .Z(n3421) );
  HS65_LS_NAND2X2 U17300 ( .A(n2596), .B(n2612), .Z(n2262) );
  HS65_LS_NAND2X2 U17301 ( .A(n1844), .B(n1860), .Z(n1510) );
  HS65_LS_NAND2X2 U17302 ( .A(n4169), .B(n4160), .Z(n3067) );
  HS65_LS_NAND2X2 U17303 ( .A(n8987), .B(n8977), .Z(n7760) );
  HS65_LS_NAND2X2 U17304 ( .A(n8938), .B(n8917), .Z(n7777) );
  HS65_LS_NAND2X2 U17305 ( .A(n8998), .B(n8987), .Z(n8136) );
  HS65_LS_NAND2X2 U17306 ( .A(n1841), .B(n1863), .Z(n1775) );
  HS65_LS_NAND2X2 U17307 ( .A(n2593), .B(n2615), .Z(n2527) );
  HS65_LS_NAND2X2 U17308 ( .A(n1468), .B(n1484), .Z(n1134) );
  HS65_LS_NAND2X2 U17309 ( .A(n2220), .B(n2236), .Z(n1886) );
  HS65_LS_NAND2X2 U17310 ( .A(n4211), .B(n4212), .Z(n3101) );
  HS65_LS_NAND2X2 U17311 ( .A(n5816), .B(n5811), .Z(n4544) );
  HS65_LS_NAND2X2 U17312 ( .A(n5934), .B(n5924), .Z(n4510) );
  HS65_LS_NAND2X2 U17313 ( .A(n7526), .B(n7516), .Z(n6103) );
  HS65_LS_NAND2X2 U17314 ( .A(n7467), .B(n7457), .Z(n6057) );
  HS65_LS_NAND2X2 U17315 ( .A(n7408), .B(n7403), .Z(n6137) );
  HS65_LS_NAND2X2 U17316 ( .A(n5875), .B(n5865), .Z(n4464) );
  HS65_LS_NAND2X2 U17317 ( .A(n5749), .B(n5762), .Z(n4676) );
  HS65_LS_NAND2X2 U17318 ( .A(n7341), .B(n7354), .Z(n6269) );
  HS65_LS_NAND2X2 U17319 ( .A(n5754), .B(n5749), .Z(n4488) );
  HS65_LS_NAND2X2 U17320 ( .A(n7346), .B(n7341), .Z(n6081) );
  HS65_LS_NAND2X2 U17321 ( .A(n4347), .B(n4340), .Z(n3391) );
  HS65_LS_NAND2X2 U17322 ( .A(n4274), .B(n4275), .Z(n2894) );
  HS65_LS_NAND2X2 U17323 ( .A(n5760), .B(n5737), .Z(n4719) );
  HS65_LS_NAND2X2 U17324 ( .A(n7352), .B(n7329), .Z(n6312) );
  HS65_LS_NAND2X2 U17325 ( .A(n4223), .B(n4229), .Z(n3100) );
  HS65_LS_NAND2X2 U17326 ( .A(n4167), .B(n4156), .Z(n3262) );
  HS65_LS_NAND2X2 U17327 ( .A(n5930), .B(n5931), .Z(n4512) );
  HS65_LS_NAND2X2 U17328 ( .A(n5871), .B(n5872), .Z(n4466) );
  HS65_LS_NAND2X2 U17329 ( .A(n7522), .B(n7523), .Z(n6105) );
  HS65_LS_NAND2X2 U17330 ( .A(n5822), .B(n5799), .Z(n4860) );
  HS65_LS_NAND2X2 U17331 ( .A(n7414), .B(n7391), .Z(n6453) );
  HS65_LS_NAND2X2 U17332 ( .A(n7463), .B(n7464), .Z(n6059) );
  HS65_LS_NAND2X2 U17333 ( .A(n5748), .B(n5749), .Z(n4721) );
  HS65_LS_NAND2X2 U17334 ( .A(n7340), .B(n7341), .Z(n6314) );
  HS65_LS_NAND2X2 U17335 ( .A(n5923), .B(n5924), .Z(n4990) );
  HS65_LS_NAND2X2 U17336 ( .A(n5864), .B(n5865), .Z(n4936) );
  HS65_LS_NAND2X2 U17337 ( .A(n5810), .B(n5811), .Z(n4861) );
  HS65_LS_NAND2X2 U17338 ( .A(n7515), .B(n7516), .Z(n6583) );
  HS65_LS_NAND2X2 U17339 ( .A(n7456), .B(n7457), .Z(n6529) );
  HS65_LS_NAND2X2 U17340 ( .A(n7402), .B(n7403), .Z(n6454) );
  HS65_LS_NAND2X2 U17341 ( .A(n1465), .B(n1487), .Z(n1399) );
  HS65_LS_NAND2X2 U17342 ( .A(n4334), .B(n4350), .Z(n3415) );
  HS65_LS_NAND2X2 U17343 ( .A(n4147), .B(n4150), .Z(n2924) );
  HS65_LS_NAND2X2 U17344 ( .A(n9111), .B(n9112), .Z(n8186) );
  HS65_LS_NAND2X2 U17345 ( .A(n9053), .B(n9054), .Z(n8154) );
  HS65_LS_NAND2X2 U17346 ( .A(n1489), .B(n1478), .Z(n1214) );
  HS65_LS_NAND2X2 U17347 ( .A(n2241), .B(n2230), .Z(n1966) );
  HS65_LS_NAND2X2 U17348 ( .A(n4219), .B(n4231), .Z(n2946) );
  HS65_LS_NAND2X2 U17349 ( .A(n2617), .B(n2606), .Z(n2342) );
  HS65_LS_NAND2X2 U17350 ( .A(n8936), .B(n8929), .Z(n7778) );
  HS65_LS_NAND2X2 U17351 ( .A(n4338), .B(n4347), .Z(n2854) );
  HS65_LS_NAND2X2 U17352 ( .A(n1865), .B(n1854), .Z(n1590) );
  HS65_LS_NAND2X2 U17353 ( .A(n9057), .B(n9058), .Z(n7634) );
  HS65_LS_NAND2X2 U17354 ( .A(n9115), .B(n9116), .Z(n7662) );
  HS65_LS_NAND2X2 U17355 ( .A(n5812), .B(n5820), .Z(n4543) );
  HS65_LS_NAND2X2 U17356 ( .A(n5932), .B(n5933), .Z(n4613) );
  HS65_LS_NAND2X2 U17357 ( .A(n7524), .B(n7525), .Z(n6206) );
  HS65_LS_NAND2X2 U17358 ( .A(n7465), .B(n7466), .Z(n6194) );
  HS65_LS_NAND2X2 U17359 ( .A(n7404), .B(n7412), .Z(n6136) );
  HS65_LS_NAND2X2 U17360 ( .A(n5873), .B(n5874), .Z(n4601) );
  HS65_LS_NAND2X2 U17361 ( .A(n8999), .B(n8977), .Z(n7872) );
  HS65_LS_NAND2X2 U17362 ( .A(n4150), .B(n4164), .Z(n3281) );
  HS65_LS_NAND2X2 U17363 ( .A(n8939), .B(n8938), .Z(n8525) );
  HS65_LS_NAND2X2 U17364 ( .A(n8997), .B(n9002), .Z(n8018) );
  HS65_LS_NAND2X2 U17365 ( .A(n8942), .B(n8934), .Z(n8060) );
  HS65_LS_NAND2X2 U17366 ( .A(n2217), .B(n2239), .Z(n2151) );
  HS65_LS_NAND2X2 U17367 ( .A(n8917), .B(n8918), .Z(n8556) );
  HS65_LS_NAND2X2 U17368 ( .A(n8977), .B(n8978), .Z(n8252) );
  HS65_LS_NAND2X2 U17369 ( .A(n1476), .B(n1467), .Z(n1129) );
  HS65_LS_NAND2X2 U17370 ( .A(n2604), .B(n2595), .Z(n2257) );
  HS65_LS_NAND2X2 U17371 ( .A(n2228), .B(n2219), .Z(n1881) );
  HS65_LS_NAND2X2 U17372 ( .A(n1852), .B(n1843), .Z(n1505) );
  HS65_LS_NAND2X2 U17373 ( .A(n7476), .B(n7454), .Z(n7136) );
  HS65_LS_NAND2X2 U17374 ( .A(n7349), .B(n7330), .Z(n7116) );
  HS65_LS_NAND2X2 U17375 ( .A(n5757), .B(n5738), .Z(n5524) );
  HS65_LS_NAND2X2 U17376 ( .A(n5943), .B(n5921), .Z(n5565) );
  HS65_LS_NAND2X2 U17377 ( .A(n7535), .B(n7513), .Z(n7157) );
  HS65_LS_NAND2X2 U17378 ( .A(n5884), .B(n5862), .Z(n5544) );
  HS65_LS_NAND2X2 U17379 ( .A(n5819), .B(n5800), .Z(n5589) );
  HS65_LS_NAND2X2 U17380 ( .A(n7411), .B(n7392), .Z(n7181) );
  HS65_LS_NAND2X2 U17381 ( .A(n2602), .B(n2603), .Z(n2286) );
  HS65_LS_NAND2X2 U17382 ( .A(n1850), .B(n1851), .Z(n1534) );
  HS65_LS_NAND2X2 U17383 ( .A(n4282), .B(n4274), .Z(n3146) );
  HS65_LS_NAND2X2 U17384 ( .A(n2618), .B(n2615), .Z(n2301) );
  HS65_LS_NAND2X2 U17385 ( .A(n1866), .B(n1863), .Z(n1549) );
  HS65_LS_NAND2X2 U17386 ( .A(n2236), .B(n2230), .Z(n1995) );
  HS65_LS_NAND2X2 U17387 ( .A(n1484), .B(n1478), .Z(n1243) );
  HS65_LS_NAND2X2 U17388 ( .A(n2612), .B(n2606), .Z(n2371) );
  HS65_LS_NAND2X2 U17389 ( .A(n1860), .B(n1854), .Z(n1619) );
  HS65_LS_NAND2X2 U17390 ( .A(n8926), .B(n8921), .Z(n7779) );
  HS65_LS_NAND2X2 U17391 ( .A(n2593), .B(n2604), .Z(n2299) );
  HS65_LS_NAND2X2 U17392 ( .A(n1841), .B(n1852), .Z(n1547) );
  HS65_LS_NAND2X2 U17393 ( .A(n8994), .B(n8981), .Z(n7762) );
  HS65_LS_NAND2X2 U17394 ( .A(n8929), .B(n8938), .Z(n7953) );
  HS65_LS_NAND2X2 U17395 ( .A(n1474), .B(n1475), .Z(n1158) );
  HS65_LS_NAND2X2 U17396 ( .A(n2226), .B(n2227), .Z(n1910) );
  HS65_LS_NAND2X2 U17397 ( .A(n1490), .B(n1487), .Z(n1173) );
  HS65_LS_NAND2X2 U17398 ( .A(n9059), .B(n9037), .Z(n7638) );
  HS65_LS_NAND2X2 U17399 ( .A(n9117), .B(n9095), .Z(n7666) );
  HS65_LS_NAND2X2 U17400 ( .A(n4290), .B(n4281), .Z(n3329) );
  HS65_LS_NAND2X2 U17401 ( .A(n9000), .B(n8987), .Z(n7870) );
  HS65_LS_NAND2X2 U17402 ( .A(n5924), .B(n5945), .Z(n5008) );
  HS65_LS_NAND2X2 U17403 ( .A(n5865), .B(n5886), .Z(n4894) );
  HS65_LS_NAND2X2 U17404 ( .A(n7516), .B(n7537), .Z(n6601) );
  HS65_LS_NAND2X2 U17405 ( .A(n7457), .B(n7478), .Z(n6487) );
  HS65_LS_NAND2X2 U17406 ( .A(n5811), .B(n5824), .Z(n4880) );
  HS65_LS_NAND2X2 U17407 ( .A(n7403), .B(n7416), .Z(n6473) );
  HS65_LS_NAND2X2 U17408 ( .A(n4169), .B(n4164), .Z(n3282) );
  HS65_LS_NAND2X2 U17409 ( .A(n4336), .B(n4337), .Z(n3007) );
  HS65_LS_NAND2X2 U17410 ( .A(n8995), .B(n8980), .Z(n8130) );
  HS65_LS_NAND2X2 U17411 ( .A(n1465), .B(n1476), .Z(n1171) );
  HS65_LS_NAND2X2 U17412 ( .A(n2603), .B(n2616), .Z(n2314) );
  HS65_LS_NAND2X2 U17413 ( .A(n1851), .B(n1864), .Z(n1562) );
  HS65_LS_NAND2X2 U17414 ( .A(n4294), .B(n4293), .Z(n3148) );
  HS65_LS_NAND2X2 U17415 ( .A(n4229), .B(n4231), .Z(n3127) );
  HS65_LS_NAND2X2 U17416 ( .A(n9030), .B(n9061), .Z(n8699) );
  HS65_LS_NAND2X2 U17417 ( .A(n9088), .B(n9119), .Z(n8787) );
  HS65_LS_NAND2X2 U17418 ( .A(n9055), .B(n9052), .Z(n7842) );
  HS65_LS_NAND2X2 U17419 ( .A(n9113), .B(n9110), .Z(n7881) );
  HS65_LS_NAND2X2 U17420 ( .A(n2242), .B(n2239), .Z(n1925) );
  HS65_LS_NAND2X2 U17421 ( .A(n4221), .B(n4213), .Z(n2877) );
  HS65_LS_NAND2X2 U17422 ( .A(n4277), .B(n4278), .Z(n2989) );
  HS65_LS_NAND2X2 U17423 ( .A(n4158), .B(n4163), .Z(n3044) );
  HS65_LS_NAND2X2 U17424 ( .A(n4353), .B(n4350), .Z(n3189) );
  HS65_LS_NAND2X2 U17425 ( .A(n9059), .B(n9056), .Z(n7847) );
  HS65_LS_NAND2X2 U17426 ( .A(n9117), .B(n9114), .Z(n7886) );
  HS65_LS_NAND2X2 U17427 ( .A(n8998), .B(n8978), .Z(n8030) );
  HS65_LS_NAND2X2 U17428 ( .A(n8997), .B(n8980), .Z(n7871) );
  HS65_LS_NAND2X2 U17429 ( .A(n4148), .B(n4164), .Z(n3057) );
  HS65_LS_NAND2X2 U17430 ( .A(n8941), .B(n8942), .Z(n7961) );
  HS65_LS_NAND2X2 U17431 ( .A(n4147), .B(n4148), .Z(n3263) );
  HS65_LS_NAND2X2 U17432 ( .A(n4169), .B(n4147), .Z(n3297) );
  HS65_LS_NAND2X2 U17433 ( .A(n2616), .B(n2617), .Z(n2263) );
  HS65_LS_NAND2X2 U17434 ( .A(n1864), .B(n1865), .Z(n1511) );
  HS65_LS_NAND2X2 U17435 ( .A(n2217), .B(n2228), .Z(n1923) );
  HS65_LS_NAND2X2 U17436 ( .A(n1475), .B(n1488), .Z(n1186) );
  HS65_LS_NAND2X2 U17437 ( .A(n2227), .B(n2240), .Z(n1938) );
  HS65_LS_NAND2X2 U17438 ( .A(n8926), .B(n8940), .Z(n8379) );
  HS65_LS_NAND2X2 U17439 ( .A(n4279), .B(n4290), .Z(n2899) );
  HS65_LS_NAND2X2 U17440 ( .A(n8936), .B(n8917), .Z(n7959) );
  HS65_LS_NAND2X2 U17441 ( .A(n8994), .B(n8995), .Z(n8315) );
  HS65_LS_NAND2X2 U17442 ( .A(n2592), .B(n2613), .Z(n2250) );
  HS65_LS_NAND2X2 U17443 ( .A(n1840), .B(n1861), .Z(n1498) );
  HS65_LS_NAND2X2 U17444 ( .A(n5750), .B(n5758), .Z(n4487) );
  HS65_LS_NAND2X2 U17445 ( .A(n7342), .B(n7350), .Z(n6080) );
  HS65_LS_NAND2X2 U17446 ( .A(n8996), .B(n8997), .Z(n7859) );
  HS65_LS_NAND2X2 U17447 ( .A(n8927), .B(n8920), .Z(n8326) );
  HS65_LS_NAND2X2 U17448 ( .A(n8940), .B(n8934), .Z(n8051) );
  HS65_LS_NAND2X2 U17449 ( .A(n9053), .B(n9057), .Z(n8159) );
  HS65_LS_NAND2X2 U17450 ( .A(n9111), .B(n9115), .Z(n8191) );
  HS65_LS_NAND2X2 U17451 ( .A(n9038), .B(n9056), .Z(n7687) );
  HS65_LS_NAND2X2 U17452 ( .A(n9096), .B(n9114), .Z(n7725) );
  HS65_LS_NAND2X2 U17453 ( .A(n5931), .B(n5921), .Z(n4783) );
  HS65_LS_NAND2X2 U17454 ( .A(n5872), .B(n5862), .Z(n4744) );
  HS65_LS_NAND2X2 U17455 ( .A(n5799), .B(n5800), .Z(n4637) );
  HS65_LS_NAND2X2 U17456 ( .A(n7523), .B(n7513), .Z(n6376) );
  HS65_LS_NAND2X2 U17457 ( .A(n7464), .B(n7454), .Z(n6337) );
  HS65_LS_NAND2X2 U17458 ( .A(n7391), .B(n7392), .Z(n6230) );
  HS65_LS_NAND2X2 U17459 ( .A(n2612), .B(n2616), .Z(n2328) );
  HS65_LS_NAND2X2 U17460 ( .A(n1860), .B(n1864), .Z(n1576) );
  HS65_LS_NAND2X2 U17461 ( .A(n1488), .B(n1489), .Z(n1135) );
  HS65_LS_NAND2X2 U17462 ( .A(n2240), .B(n2241), .Z(n1887) );
  HS65_LS_NAND2X2 U17463 ( .A(n5737), .B(n5738), .Z(n4559) );
  HS65_LS_NAND2X2 U17464 ( .A(n7329), .B(n7330), .Z(n6152) );
  HS65_LS_NAND2X2 U17465 ( .A(n1464), .B(n1485), .Z(n1122) );
  HS65_LS_NAND2X2 U17466 ( .A(n2216), .B(n2237), .Z(n1874) );
  HS65_LS_NAND2X2 U17467 ( .A(n8996), .B(n9001), .Z(n8663) );
  HS65_LS_NAND2X2 U17468 ( .A(n9050), .B(n9051), .Z(n7645) );
  HS65_LS_NAND2X2 U17469 ( .A(n9108), .B(n9109), .Z(n7673) );
  HS65_LS_NAND2X2 U17470 ( .A(n4335), .B(n4334), .Z(n3893) );
  HS65_LS_NAND2X2 U17471 ( .A(n1465), .B(n1486), .Z(n1156) );
  HS65_LS_NAND2X2 U17472 ( .A(n2593), .B(n2614), .Z(n2284) );
  HS65_LS_NAND2X2 U17473 ( .A(n2217), .B(n2238), .Z(n1908) );
  HS65_LS_NAND2X2 U17474 ( .A(n1841), .B(n1862), .Z(n1532) );
  HS65_LS_NAND2X2 U17475 ( .A(n9110), .B(n9117), .Z(n8181) );
  HS65_LS_NAND2X2 U17476 ( .A(n9052), .B(n9059), .Z(n8149) );
  HS65_LS_NAND2X2 U17477 ( .A(n9052), .B(n9038), .Z(n7833) );
  HS65_LS_NAND2X2 U17478 ( .A(n9110), .B(n9096), .Z(n7932) );
  HS65_LS_NAND2X2 U17479 ( .A(n1484), .B(n1488), .Z(n1200) );
  HS65_LS_NAND2X2 U17480 ( .A(n2236), .B(n2240), .Z(n1952) );
  HS65_LS_NAND2X2 U17481 ( .A(n4156), .B(n4165), .Z(n3066) );
  HS65_LS_NAND2X2 U17482 ( .A(n8995), .B(n9002), .Z(n8119) );
  HS65_LS_NAND2X2 U17483 ( .A(n4351), .B(n4352), .Z(n2855) );
  HS65_LS_NAND2X2 U17484 ( .A(n4287), .B(n4288), .Z(n2900) );
  HS65_LS_NAND2X2 U17485 ( .A(n4230), .B(n4228), .Z(n3905) );
  HS65_LS_NAND2X2 U17486 ( .A(n7479), .B(n7456), .Z(n6063) );
  HS65_LS_NAND2X2 U17487 ( .A(n5751), .B(n5748), .Z(n4495) );
  HS65_LS_NAND2X2 U17488 ( .A(n5946), .B(n5923), .Z(n4516) );
  HS65_LS_NAND2X2 U17489 ( .A(n7538), .B(n7515), .Z(n6109) );
  HS65_LS_NAND2X2 U17490 ( .A(n5887), .B(n5864), .Z(n4470) );
  HS65_LS_NAND2X2 U17491 ( .A(n7343), .B(n7340), .Z(n6088) );
  HS65_LS_NAND2X2 U17492 ( .A(n5813), .B(n5810), .Z(n4535) );
  HS65_LS_NAND2X2 U17493 ( .A(n7405), .B(n7402), .Z(n6128) );
  HS65_LS_NAND2X2 U17494 ( .A(n4335), .B(n4348), .Z(n2842) );
  HS65_LS_NAND2X2 U17495 ( .A(n4163), .B(n4165), .Z(n3053) );
  HS65_LS_NAND2X2 U17496 ( .A(n4338), .B(n4339), .Z(n2850) );
  HS65_LS_NAND2X2 U17497 ( .A(n5753), .B(n5761), .Z(n4722) );
  HS65_LS_NAND2X2 U17498 ( .A(n7345), .B(n7353), .Z(n6315) );
  HS65_LS_NAND2X2 U17499 ( .A(n5757), .B(n5753), .Z(n4561) );
  HS65_LS_NAND2X2 U17500 ( .A(n7349), .B(n7345), .Z(n6154) );
  HS65_LS_NAND2X2 U17501 ( .A(n8988), .B(n8999), .Z(n8267) );
  HS65_LS_NAND2X2 U17502 ( .A(n8989), .B(n8977), .Z(n7857) );
  HS65_LS_NAND2X2 U17503 ( .A(n4347), .B(n4351), .Z(n3208) );
  HS65_LS_NAND2X2 U17504 ( .A(n9116), .B(n9088), .Z(n7660) );
  HS65_LS_NAND2X2 U17505 ( .A(n9058), .B(n9030), .Z(n7632) );
  HS65_LS_NAND2X2 U17506 ( .A(n9029), .B(n9044), .Z(n7642) );
  HS65_LS_NAND2X2 U17507 ( .A(n9087), .B(n9102), .Z(n7670) );
  HS65_LS_NAND2X2 U17508 ( .A(n4213), .B(n4230), .Z(n3538) );
  HS65_LS_NAND2X2 U17509 ( .A(n4278), .B(n4287), .Z(n3778) );
  HS65_LS_NAND2X2 U17510 ( .A(n8939), .B(n8928), .Z(n8571) );
  HS65_LS_NAND2X2 U17511 ( .A(n4276), .B(n4291), .Z(n2887) );
  HS65_LS_NAND2X2 U17512 ( .A(n4336), .B(n4339), .Z(n3845) );
  HS65_LS_NAND2X2 U17513 ( .A(n7346), .B(n7350), .Z(n6634) );
  HS65_LS_NAND2X2 U17514 ( .A(n5754), .B(n5758), .Z(n5041) );
  HS65_LS_NAND2X2 U17515 ( .A(n8935), .B(n8918), .Z(n8069) );
  HS65_LS_NAND2X2 U17516 ( .A(n7467), .B(n7466), .Z(n6872) );
  HS65_LS_NAND2X2 U17517 ( .A(n5934), .B(n5933), .Z(n5395) );
  HS65_LS_NAND2X2 U17518 ( .A(n7408), .B(n7412), .Z(n6755) );
  HS65_LS_NAND2X2 U17519 ( .A(n5816), .B(n5820), .Z(n5163) );
  HS65_LS_NAND2X2 U17520 ( .A(n7526), .B(n7525), .Z(n6987) );
  HS65_LS_NAND2X2 U17521 ( .A(n5875), .B(n5874), .Z(n5280) );
  HS65_LS_NAND2X2 U17522 ( .A(n4225), .B(n4223), .Z(n2944) );
  HS65_LS_NAND2X2 U17523 ( .A(n4341), .B(n4333), .Z(n3187) );
  HS65_LSS_XOR2X3 U17524 ( .A(n936), .B(n1098), .Z(n1050) );
  HS65_LSS_XOR2X3 U17525 ( .A(n935), .B(n1107), .Z(n1068) );
  HS65_LSS_XOR2X3 U17526 ( .A(n940), .B(n1093), .Z(n1040) );
  HS65_LS_NAND2X2 U17527 ( .A(n8989), .B(n9000), .Z(n7761) );
  HS65_LS_NAND2X2 U17528 ( .A(n8980), .B(n8981), .Z(n8019) );
  HS65_LS_NAND2X2 U17529 ( .A(n8920), .B(n8921), .Z(n8061) );
  HS65_LS_NAND2X2 U17530 ( .A(n5930), .B(n5940), .Z(n5626) );
  HS65_LS_NAND2X2 U17531 ( .A(n5871), .B(n5881), .Z(n5599) );
  HS65_LS_NAND2X2 U17532 ( .A(n5822), .B(n5823), .Z(n5582) );
  HS65_LS_NAND2X2 U17533 ( .A(n7522), .B(n7532), .Z(n7218) );
  HS65_LS_NAND2X2 U17534 ( .A(n7463), .B(n7473), .Z(n7191) );
  HS65_LS_NAND2X2 U17535 ( .A(n7414), .B(n7415), .Z(n7174) );
  HS65_LSS_XOR2X3 U17536 ( .A(n958), .B(n1807), .Z(n1002) );
  HS65_LS_NAND4ABX3 U17537 ( .A(n1808), .B(n1809), .C(n1810), .D(n1811), .Z(
        n1807) );
  HS65_LS_NOR4ABX2 U17538 ( .A(n1552), .B(n1687), .C(n1812), .D(n1701), .Z(
        n1811) );
  HS65_LS_MX41X4 U17539 ( .D0(n825), .S0(n842), .D1(n826), .S1(n834), .D2(n845), .S2(n818), .D3(n846), .S3(n1554), .Z(n1809) );
  HS65_LS_NAND2X2 U17540 ( .A(n9044), .B(n9061), .Z(n7697) );
  HS65_LS_NAND2X2 U17541 ( .A(n9102), .B(n9119), .Z(n7735) );
  HS65_LS_NAND2X2 U17542 ( .A(n4276), .B(n4275), .Z(n3776) );
  HS65_LSS_XOR2X3 U17543 ( .A(n941), .B(n1088), .Z(n1030) );
  HS65_LSS_XOR2X3 U17544 ( .A(n943), .B(n1084), .Z(n1022) );
  HS65_LS_NAND2X2 U17545 ( .A(n5939), .B(n5940), .Z(n4503) );
  HS65_LS_NAND2X2 U17546 ( .A(n5880), .B(n5881), .Z(n4457) );
  HS65_LS_NAND2X2 U17547 ( .A(n7531), .B(n7532), .Z(n6096) );
  HS65_LS_NAND2X2 U17548 ( .A(n7472), .B(n7473), .Z(n6050) );
  HS65_LS_NAND2X2 U17549 ( .A(n5818), .B(n5823), .Z(n4835) );
  HS65_LS_NAND2X2 U17550 ( .A(n7410), .B(n7415), .Z(n6428) );
  HS65_LSS_XOR2X3 U17551 ( .A(n942), .B(n1087), .Z(n1028) );
  HS65_LSS_XOR2X3 U17552 ( .A(n937), .B(n1097), .Z(n1048) );
  HS65_LSS_XOR2X3 U17553 ( .A(n939), .B(n1095), .Z(n1044) );
  HS65_LSS_XOR2X3 U17554 ( .A(n957), .B(n1867), .Z(n1003) );
  HS65_LS_NAND4ABX3 U17555 ( .A(n1868), .B(n1869), .C(n1870), .D(n1871), .Z(
        n1867) );
  HS65_LS_NAND4ABX3 U17556 ( .A(n1889), .B(n1890), .C(n1891), .D(n1892), .Z(
        n1868) );
  HS65_LS_OAI212X3 U17557 ( .A(n1879), .B(n1880), .C(n1881), .D(n1882), .E(
        n1883), .Z(n1869) );
  HS65_LSS_XOR2X3 U17558 ( .A(n959), .B(n1782), .Z(n1001) );
  HS65_LS_NAND4ABX3 U17559 ( .A(n1783), .B(n1784), .C(n1785), .D(n1786), .Z(
        n1782) );
  HS65_LS_AOI222X2 U17560 ( .A(n836), .B(n814), .C(n833), .D(n1805), .E(n845), 
        .F(n813), .Z(n1785) );
  HS65_LS_CB4I6X4 U17561 ( .A(n817), .B(n822), .C(n844), .D(n1703), .Z(n1783)
         );
  HS65_LSS_XOR2X3 U17562 ( .A(n952), .B(n2534), .Z(n1017) );
  HS65_LS_NAND4ABX3 U17563 ( .A(n2535), .B(n2536), .C(n2537), .D(n2538), .Z(
        n2534) );
  HS65_LS_AOI222X2 U17564 ( .A(n918), .B(n896), .C(n915), .D(n2557), .E(n927), 
        .F(n895), .Z(n2537) );
  HS65_LS_CB4I6X4 U17565 ( .A(n899), .B(n904), .C(n926), .D(n2455), .Z(n2535)
         );
  HS65_LS_NAND2X2 U17566 ( .A(n4157), .B(n4155), .Z(n2925) );
  HS65_LSS_XOR2X3 U17567 ( .A(n938), .B(n1096), .Z(n1046) );
  HS65_LS_NAND2X2 U17568 ( .A(n9112), .B(n9087), .Z(n7885) );
  HS65_LS_NAND2X2 U17569 ( .A(n9054), .B(n9029), .Z(n7846) );
  HS65_LS_NAND2X2 U17570 ( .A(n1474), .B(n1469), .Z(n1312) );
  HS65_LS_NAND2X2 U17571 ( .A(n2226), .B(n2221), .Z(n2064) );
  HS65_LS_NAND2X2 U17572 ( .A(n2602), .B(n2597), .Z(n2440) );
  HS65_LS_NAND2X2 U17573 ( .A(n1850), .B(n1845), .Z(n1688) );
  HS65_LS_NAND2X2 U17574 ( .A(n5943), .B(n5941), .Z(n4784) );
  HS65_LS_NAND2X2 U17575 ( .A(n5884), .B(n5882), .Z(n4745) );
  HS65_LS_NAND2X2 U17576 ( .A(n5819), .B(n5815), .Z(n4638) );
  HS65_LS_NAND2X2 U17577 ( .A(n7535), .B(n7533), .Z(n6377) );
  HS65_LS_NAND2X2 U17578 ( .A(n7476), .B(n7474), .Z(n6338) );
  HS65_LS_NAND2X2 U17579 ( .A(n7411), .B(n7407), .Z(n6231) );
  HS65_LSS_XOR2X3 U17580 ( .A(n956), .B(n1894), .Z(n1004) );
  HS65_LS_NAND4ABX3 U17581 ( .A(n1895), .B(n1896), .C(n1897), .D(n1898), .Z(
        n1894) );
  HS65_LS_CBI4I1X3 U17582 ( .A(n1910), .B(n1880), .C(n1911), .D(n1912), .Z(
        n1895) );
  HS65_LS_AOI212X2 U17583 ( .A(n805), .B(n771), .C(n802), .D(n783), .E(n1904), 
        .Z(n1897) );
  HS65_LS_NAND2X2 U17584 ( .A(n4221), .B(n4222), .Z(n3486) );
  HS65_LS_NAND2X2 U17585 ( .A(n4274), .B(n4291), .Z(n3174) );
  HS65_LS_NAND2X2 U17586 ( .A(n4226), .B(n4224), .Z(n3123) );
  HS65_LS_NAND2X2 U17587 ( .A(n4277), .B(n4280), .Z(n3728) );
  HS65_LS_NAND2X2 U17588 ( .A(n4282), .B(n4292), .Z(n2987) );
  HS65_LS_NAND2X2 U17589 ( .A(n4225), .B(n4220), .Z(n2875) );
  HS65_LS_NAND2X2 U17590 ( .A(n4341), .B(n4349), .Z(n3005) );
  HS65_LS_NOR2X2 U17591 ( .A(n183), .B(n178), .Z(n4168) );
  HS65_LSS_XOR2X3 U17592 ( .A(n2134), .B(n955), .Z(n1008) );
  HS65_LS_NOR4ABX2 U17593 ( .A(n2135), .B(n2136), .C(n2137), .D(n2138), .Z(
        n2134) );
  HS65_LS_CBI4I1X3 U17594 ( .A(n1953), .B(n1881), .C(n1907), .D(n2086), .Z(
        n2138) );
  HS65_LS_CBI4I6X2 U17595 ( .A(n778), .B(n2108), .C(n799), .D(n2157), .Z(n2135) );
  HS65_LSS_XOR2X3 U17596 ( .A(n1537), .B(n962), .Z(n997) );
  HS65_LS_NOR3X1 U17597 ( .A(n1538), .B(n1539), .C(n1540), .Z(n1537) );
  HS65_LS_NAND4ABX3 U17598 ( .A(n1565), .B(n1566), .C(n1567), .D(n1568), .Z(
        n1538) );
  HS65_LS_OAI212X3 U17599 ( .A(n1505), .B(n1510), .C(n1532), .D(n1562), .E(
        n1563), .Z(n1539) );
  HS65_LSS_XOR2X3 U17600 ( .A(n1758), .B(n960), .Z(n1000) );
  HS65_LS_NOR4ABX2 U17601 ( .A(n1759), .B(n1760), .C(n1761), .D(n1762), .Z(
        n1758) );
  HS65_LS_CBI4I1X3 U17602 ( .A(n1577), .B(n1505), .C(n1531), .D(n1710), .Z(
        n1762) );
  HS65_LS_CBI4I6X2 U17603 ( .A(n819), .B(n1732), .C(n840), .D(n1781), .Z(n1759) );
  HS65_LSS_XNOR2X3 U17604 ( .A(n997), .B(n945), .Z(n1093) );
  HS65_LSS_XNOR2X3 U17605 ( .A(n1000), .B(n944), .Z(n1096) );
  HS65_LSS_XNOR2X3 U17606 ( .A(n992), .B(n947), .Z(n1088) );
  HS65_LSS_XNOR2X3 U17607 ( .A(n989), .B(n949), .Z(n1085) );
  HS65_LSS_XNOR2X3 U17608 ( .A(n990), .B(n948), .Z(n1086) );
  HS65_LSS_XOR2X3 U17609 ( .A(n961), .B(n1641), .Z(n999) );
  HS65_LS_NAND4ABX3 U17610 ( .A(n1642), .B(n1643), .C(n1644), .D(n1645), .Z(
        n1641) );
  HS65_LS_MX41X4 U17611 ( .D0(n815), .S0(n839), .D1(n843), .S1(n827), .D2(n813), .S2(n834), .D3(n845), .S3(n1554), .Z(n1643) );
  HS65_LS_AOI212X2 U17612 ( .A(n828), .B(n1646), .C(n844), .D(n1623), .E(n1647), .Z(n1645) );
  HS65_LSS_XOR2X3 U17613 ( .A(n2674), .B(n790), .Z(n9843) );
  HS65_LS_NOR3AX2 U17614 ( .A(n981), .B(n978), .C(n974), .Z(n984) );
  HS65_LS_NAND2X2 U17615 ( .A(n981), .B(n974), .Z(n982) );
  HS65_LS_NAND2X2 U17616 ( .A(\u0/r0/rcnt [2]), .B(n974), .Z(n977) );
  HS65_LS_OAI311X2 U17617 ( .A(n982), .B(n972), .C(n978), .D(n983), .E(n9859), 
        .Z(\u0/rcon [24]) );
  HS65_LS_NAND2X2 U17618 ( .A(n978), .B(n9860), .Z(n975) );
  HS65_LS_NAND3X2 U17619 ( .A(n9865), .B(n972), .C(n984), .Z(n979) );
  HS65_LS_NOR2X6 U17620 ( .A(n5), .B(n2619), .Z(n2621) );
  HS65_LS_OAI13X1 U17621 ( .A(n976), .B(n982), .C(n978), .D(n980), .Z(
        \u0/rcon [25]) );
  HS65_LS_NAND2X2 U17622 ( .A(n9859), .B(n972), .Z(n976) );
  HS65_LS_OAI13X1 U17623 ( .A(n978), .B(n972), .C(n977), .D(n980), .Z(
        \u0/rcon [28]) );
  HS65_LS_OAI13X1 U17624 ( .A(n975), .B(n972), .C(n982), .D(n979), .Z(
        \u0/rcon [26]) );
  HS65_LS_IVX2 U17625 ( .A(n978), .Z(n971) );
  HS65_LS_NOR3X1 U17626 ( .A(n977), .B(n971), .C(n972), .Z(\u0/rcon [30]) );
  HS65_LS_IVX9 U17627 ( .A(n2619), .Z(n2) );
  HS65_LS_IVX2 U17628 ( .A(n2623), .Z(n3) );
  HS65_LS_NOR2X2 U17629 ( .A(n981), .B(n9846), .Z(\u0/r0/rcnt [2]) );
  HS65_LS_OA12X4 U17630 ( .A(n9858), .B(n983), .C(n979), .Z(n980) );
  HS65_LS_NOR2X2 U17631 ( .A(n9846), .B(n974), .Z(\u0/r0/rcnt [3]) );
  HS65_LS_BFX4 U17632 ( .A(n9148), .Z(n9146) );
  HS65_LS_NOR2X2 U17633 ( .A(n9382), .B(n9373), .Z(n8977) );
  HS65_LS_NOR2X2 U17634 ( .A(n9403), .B(sa02[6]), .Z(n8917) );
  HS65_LS_NOR2X2 U17635 ( .A(n339), .B(n9356), .Z(n8938) );
  HS65_LS_NOR2X2 U17636 ( .A(n9375), .B(n9348), .Z(n8989) );
  HS65_LS_NOR2X2 U17637 ( .A(n9357), .B(n9356), .Z(n8936) );
  HS65_LS_NOR2X2 U17638 ( .A(n933), .B(n9183), .Z(n2616) );
  HS65_LS_NOR2X2 U17639 ( .A(n851), .B(n9338), .Z(n1864) );
  HS65_LS_NOR2X2 U17640 ( .A(n931), .B(n9181), .Z(n2612) );
  HS65_LS_NOR2X2 U17641 ( .A(n849), .B(n9339), .Z(n1860) );
  HS65_LS_NOR2X2 U17642 ( .A(n850), .B(n9185), .Z(n1865) );
  HS65_LS_NOR2X2 U17643 ( .A(n932), .B(n9179), .Z(n2617) );
  HS65_LS_NOR2X2 U17644 ( .A(n9181), .B(n9179), .Z(n2603) );
  HS65_LS_NOR2X2 U17645 ( .A(n9339), .B(n9185), .Z(n1851) );
  HS65_LS_NOR2X2 U17646 ( .A(n9401), .B(n9376), .Z(n8980) );
  HS65_LS_NOR2X2 U17647 ( .A(n163), .B(n9310), .Z(n4169) );
  HS65_LS_NOR2X2 U17648 ( .A(n384), .B(n9348), .Z(n8987) );
  HS65_LS_NOR2X2 U17649 ( .A(n891), .B(n9175), .Z(n1489) );
  HS65_LS_NOR2X2 U17650 ( .A(n809), .B(n9186), .Z(n2241) );
  HS65_LS_NOR2X2 U17651 ( .A(n9172), .B(n9175), .Z(n1475) );
  HS65_LS_NOR2X2 U17652 ( .A(n9393), .B(n9186), .Z(n2227) );
  HS65_LS_NOR2X2 U17653 ( .A(n892), .B(n9386), .Z(n1488) );
  HS65_LS_NOR2X2 U17654 ( .A(n810), .B(n9171), .Z(n2240) );
  HS65_LS_NOR2X2 U17655 ( .A(n890), .B(n9172), .Z(n1484) );
  HS65_LS_NOR2X2 U17656 ( .A(n808), .B(n9393), .Z(n2236) );
  HS65_LS_NOR2X2 U17657 ( .A(n604), .B(n9347), .Z(n9054) );
  HS65_LS_NOR2X2 U17658 ( .A(n117), .B(n9245), .Z(n9112) );
  HS65_LS_NOR2X2 U17659 ( .A(n621), .B(n9322), .Z(n9052) );
  HS65_LS_NOR2X2 U17660 ( .A(n134), .B(sa13[2]), .Z(n9110) );
  HS65_LS_NOR2X2 U17661 ( .A(n9343), .B(n9365), .Z(n4338) );
  HS65_LS_NOR2X2 U17662 ( .A(n333), .B(sa02[6]), .Z(n8939) );
  HS65_LS_NOR2X2 U17663 ( .A(n9341), .B(n9358), .Z(n4350) );
  HS65_LS_NOR2X2 U17664 ( .A(n9361), .B(n9377), .Z(n4231) );
  HS65_LS_NOR2X2 U17665 ( .A(n9336), .B(n9243), .Z(n8920) );
  HS65_LS_NOR2X2 U17666 ( .A(n162), .B(n9299), .Z(n4164) );
  HS65_LS_NOR2X2 U17667 ( .A(n9314), .B(n9313), .Z(n9116) );
  HS65_LS_NOR2X2 U17668 ( .A(n9246), .B(n9329), .Z(n9058) );
  HS65_LS_NOR2X2 U17669 ( .A(n208), .B(n9366), .Z(n4228) );
  HS65_LS_NOR2X2 U17670 ( .A(n428), .B(n9355), .Z(n4352) );
  HS65_LS_NOR2X2 U17671 ( .A(n652), .B(n9340), .Z(n4288) );
  HS65_LS_NOR2X2 U17672 ( .A(sa03[3]), .B(sa03[2]), .Z(n4163) );
  HS65_LS_NOR2X2 U17673 ( .A(n449), .B(n9378), .Z(n4334) );
  HS65_LS_NOR2X2 U17674 ( .A(n672), .B(n9324), .Z(n4274) );
  HS65_LS_NOR2X2 U17675 ( .A(n9323), .B(n9340), .Z(n4278) );
  HS65_LS_NOR2X2 U17676 ( .A(n405), .B(n9371), .Z(n8995) );
  HS65_LS_NOR2X2 U17677 ( .A(n9387), .B(n9366), .Z(n4213) );
  HS65_LS_NOR2X2 U17678 ( .A(n361), .B(n9344), .Z(n8940) );
  HS65_LS_NOR2X2 U17679 ( .A(n429), .B(n9359), .Z(n4347) );
  HS65_LS_NOR2X2 U17680 ( .A(n934), .B(n9170), .Z(n2602) );
  HS65_LS_NOR2X2 U17681 ( .A(n9183), .B(n9170), .Z(n2596) );
  HS65_LS_NOR2X2 U17682 ( .A(n9177), .B(n9184), .Z(n1863) );
  HS65_LS_NOR2X2 U17683 ( .A(n9166), .B(n9169), .Z(n2615) );
  HS65_LS_NOR2X2 U17684 ( .A(n914), .B(n9169), .Z(n2604) );
  HS65_LS_NOR2X2 U17685 ( .A(n832), .B(n9184), .Z(n1852) );
  HS65_LS_NOR2X2 U17686 ( .A(n338), .B(n9403), .Z(n8929) );
  HS65_LS_OAI22X1 U17687 ( .A(n7539), .B(n9146), .C(n9137), .D(n7540), .Z(
        sa02[7]) );
  HS65_LSS_XNOR2X3 U17688 ( .A(n9283), .B(n9652), .Z(n7539) );
  HS65_LSS_XNOR3X2 U17689 ( .A(n3014), .B(n7541), .C(n7542), .Z(n7540) );
  HS65_LSS_XOR3X2 U17690 ( .A(n2815), .B(n9283), .C(n2816), .Z(n7541) );
  HS65_LS_OAI22X1 U17691 ( .A(n4354), .B(n9143), .C(n9139), .D(n4355), .Z(
        sa00[7]) );
  HS65_LSS_XOR2X3 U17692 ( .A(n970), .B(n9716), .Z(n4354) );
  HS65_LSS_XNOR3X2 U17693 ( .A(n3543), .B(n4356), .C(n4357), .Z(n4355) );
  HS65_LSS_XOR3X2 U17694 ( .A(n2831), .B(n9248), .C(n452), .Z(n4356) );
  HS65_LS_OAI22X1 U17695 ( .A(n9570), .B(n9575), .C(n9584), .D(n9424), .Z(
        sa01[7]) );
  HS65_LSS_XOR2X3 U17696 ( .A(n951), .B(n9684), .Z(n5947) );
  HS65_LSS_XNOR3X2 U17697 ( .A(n3218), .B(n5949), .C(n5950), .Z(n5948) );
  HS65_LS_IVX2 U17698 ( .A(n9205), .Z(n951) );
  HS65_LS_NOR2X2 U17699 ( .A(n893), .B(n9394), .Z(n1474) );
  HS65_LS_NOR2X2 U17700 ( .A(n811), .B(n9188), .Z(n2226) );
  HS65_LS_NOR2X2 U17701 ( .A(n852), .B(n9182), .Z(n1850) );
  HS65_LS_NOR2X2 U17702 ( .A(n9386), .B(n9394), .Z(n1468) );
  HS65_LS_NOR2X2 U17703 ( .A(n9171), .B(n9188), .Z(n2220) );
  HS65_LS_NOR2X2 U17704 ( .A(n9338), .B(n9182), .Z(n1844) );
  HS65_LS_NOR2X2 U17705 ( .A(n9168), .B(n9174), .Z(n1487) );
  HS65_LS_NOR2X2 U17706 ( .A(n873), .B(n9174), .Z(n1476) );
  HS65_LS_IVX2 U17707 ( .A(n9190), .Z(n790) );
  HS65_LS_OAI22X1 U17708 ( .A(n6721), .B(n9145), .C(n9136), .D(n6722), .Z(
        sa31[3]) );
  HS65_LSS_XNOR2X3 U17709 ( .A(n9222), .B(n9656), .Z(n6721) );
  HS65_LSS_XNOR3X2 U17710 ( .A(n6004), .B(n6723), .C(n6406), .Z(n6722) );
  HS65_LSS_XNOR3X2 U17711 ( .A(n9222), .B(n5967), .C(n3019), .Z(n6723) );
  HS65_LS_OAI22X1 U17712 ( .A(n4362), .B(n9143), .C(n9588), .D(n4363), .Z(
        sa00[5]) );
  HS65_LSS_XOR2X3 U17713 ( .A(n968), .B(n9714), .Z(n4362) );
  HS65_LSS_XNOR3X2 U17714 ( .A(n3224), .B(n4364), .C(n4365), .Z(n4363) );
  HS65_LSS_XOR3X2 U17715 ( .A(n2782), .B(n9194), .C(n2829), .Z(n4364) );
  HS65_LS_NOR2X2 U17716 ( .A(n9383), .B(n9388), .Z(n4279) );
  HS65_LS_NOR2X2 U17717 ( .A(n382), .B(n9373), .Z(n8988) );
  HS65_LS_NOR2X2 U17718 ( .A(n206), .B(n9368), .Z(n4221) );
  HS65_LS_NOR2X2 U17719 ( .A(n418), .B(n9365), .Z(n4336) );
  HS65_LS_NOR2X2 U17720 ( .A(n642), .B(n9388), .Z(n4277) );
  HS65_LS_NOR2X2 U17721 ( .A(n605), .B(n9399), .Z(n9057) );
  HS65_LS_NOR2X2 U17722 ( .A(n118), .B(n9309), .Z(n9115) );
  HS65_LS_NOR2AX3 U17723 ( .A(n9349), .B(n9380), .Z(n5930) );
  HS65_LS_NOR2AX3 U17724 ( .A(n9351), .B(n9379), .Z(n5871) );
  HS65_LS_NOR2AX3 U17725 ( .A(n9239), .B(n9318), .Z(n7522) );
  HS65_LS_NOR2AX3 U17726 ( .A(sa23[1]), .B(n9301), .Z(n7463) );
  HS65_LS_NOR2AX3 U17727 ( .A(n9333), .B(n9312), .Z(n5822) );
  HS65_LS_NOR2AX3 U17728 ( .A(n9332), .B(n9392), .Z(n7414) );
  HS65_LS_OAI22X1 U17729 ( .A(n9569), .B(n9580), .C(n9587), .D(n9423), .Z(
        sa23[2]) );
  HS65_LSS_XOR2X3 U17730 ( .A(n831), .B(n9599), .Z(n2750) );
  HS65_LSS_XNOR3X2 U17731 ( .A(n2722), .B(n2752), .C(n2715), .Z(n2751) );
  HS65_LSS_XOR3X2 U17732 ( .A(n2667), .B(n9184), .C(n2681), .Z(n2752) );
  HS65_LS_NOR2AX3 U17733 ( .A(n9243), .B(n9336), .Z(n8941) );
  HS65_LS_NOR2AX3 U17734 ( .A(n9376), .B(n9401), .Z(n8996) );
  HS65_LS_NOR2X2 U17735 ( .A(n9180), .B(n9190), .Z(n2239) );
  HS65_LS_NOR2X2 U17736 ( .A(n9327), .B(n9324), .Z(n4293) );
  HS65_LS_NOR2X2 U17737 ( .A(n9344), .B(n9370), .Z(n8921) );
  HS65_LS_NOR2X2 U17738 ( .A(n9360), .B(n9371), .Z(n8981) );
  HS65_LS_NOR2X2 U17739 ( .A(n791), .B(n9190), .Z(n2228) );
  HS65_LS_NOR2X2 U17740 ( .A(n9359), .B(n9355), .Z(n4337) );
  HS65_LS_NOR2X2 U17741 ( .A(n9315), .B(n9310), .Z(n4150) );
  HS65_LS_OAI22X1 U17742 ( .A(n4428), .B(n9146), .C(n9139), .D(n4429), .Z(
        sa20[5]) );
  HS65_LSS_XNOR2X3 U17743 ( .A(n9215), .B(n9698), .Z(n4428) );
  HS65_LSS_XNOR3X2 U17744 ( .A(n2830), .B(n4430), .C(n4398), .Z(n4429) );
  HS65_LSS_XOR3X2 U17745 ( .A(n2781), .B(n9215), .C(n2805), .Z(n4430) );
  HS65_LS_OAI22X1 U17746 ( .A(n2737), .B(n9144), .C(n9140), .D(n2738), .Z(
        sa23[5]) );
  HS65_LSS_XOR2X3 U17747 ( .A(n850), .B(n9602), .Z(n2737) );
  HS65_LSS_XNOR3X2 U17748 ( .A(n2707), .B(n2739), .C(n2699), .Z(n2738) );
  HS65_LSS_XOR3X2 U17749 ( .A(n2647), .B(n9339), .C(n2740), .Z(n2739) );
  HS65_LS_NOR2X2 U17750 ( .A(n674), .B(n9330), .Z(n4275) );
  HS65_LS_NOR2X2 U17751 ( .A(n224), .B(n9377), .Z(n4223) );
  HS65_LS_NOR2X2 U17752 ( .A(n448), .B(n9358), .Z(n4333) );
  HS65_LS_NOR2X2 U17753 ( .A(n9307), .B(n9300), .Z(n5753) );
  HS65_LS_NOR2X2 U17754 ( .A(n9242), .B(n9372), .Z(n7345) );
  HS65_LS_NOR2X2 U17755 ( .A(n653), .B(n9323), .Z(n4290) );
  HS65_LS_NOR2X2 U17756 ( .A(n164), .B(n9315), .Z(n4148) );
  HS65_LS_NOR2X2 U17757 ( .A(n116), .B(n9314), .Z(n9087) );
  HS65_LS_NOR2X2 U17758 ( .A(n603), .B(n9246), .Z(n9029) );
  HS65_LS_NOR2X2 U17759 ( .A(n383), .B(n9382), .Z(n9000) );
  HS65_LS_OAI22X1 U17760 ( .A(n4376), .B(n9143), .C(n9138), .D(n4377), .Z(
        sa00[2]) );
  HS65_LSS_XOR2X3 U17761 ( .A(n965), .B(n9711), .Z(n4376) );
  HS65_LSS_XNOR3X2 U17762 ( .A(n3221), .B(n4378), .C(n4379), .Z(n4377) );
  HS65_LSS_XOR3X2 U17763 ( .A(n2779), .B(n9192), .C(n2826), .Z(n4378) );
  HS65_LS_OAI22X1 U17764 ( .A(n5969), .B(n9145), .C(n9137), .D(n5970), .Z(
        sa01[2]) );
  HS65_LSS_XOR2X3 U17765 ( .A(n947), .B(n9679), .Z(n5969) );
  HS65_LSS_XNOR3X2 U17766 ( .A(n3017), .B(n5971), .C(n5972), .Z(n5970) );
  HS65_LSS_XOR3X2 U17767 ( .A(n2771), .B(n9198), .C(n2818), .Z(n5971) );
  HS65_LS_NOR2AX3 U17768 ( .A(n9305), .B(n9308), .Z(n7466) );
  HS65_LS_NOR2AX3 U17769 ( .A(n9385), .B(n9389), .Z(n5933) );
  HS65_LS_NOR2AX3 U17770 ( .A(n9381), .B(n9374), .Z(n7350) );
  HS65_LS_NOR2AX3 U17771 ( .A(n9302), .B(n9319), .Z(n5758) );
  HS65_LS_NOR2AX3 U17772 ( .A(n9402), .B(n9236), .Z(n5820) );
  HS65_LS_NOR2AX3 U17773 ( .A(n9390), .B(sa12[6]), .Z(n7525) );
  HS65_LS_NOR2AX3 U17774 ( .A(sa22[7]), .B(sa22[6]), .Z(n5874) );
  HS65_LS_NOR2AX3 U17775 ( .A(sa01[7]), .B(n9235), .Z(n7412) );
  HS65_LS_NOR2X2 U17776 ( .A(n28), .B(n9311), .Z(n5748) );
  HS65_LS_NOR2X2 U17777 ( .A(n554), .B(n9367), .Z(n7340) );
  HS65_LS_NOR2X2 U17778 ( .A(n470), .B(n9326), .Z(n5923) );
  HS65_LS_NOR2X2 U17779 ( .A(n251), .B(n9364), .Z(n5864) );
  HS65_LS_NOR2X2 U17780 ( .A(n692), .B(n9400), .Z(n5810) );
  HS65_LS_NOR2X2 U17781 ( .A(n293), .B(n9335), .Z(n7515) );
  HS65_LS_NOR2X2 U17782 ( .A(n72), .B(n9398), .Z(n7456) );
  HS65_LS_NOR2X2 U17783 ( .A(n510), .B(n9395), .Z(n7402) );
  HS65_LS_OAI22X1 U17784 ( .A(n5955), .B(n9146), .C(n9137), .D(n5956), .Z(
        sa01[5]) );
  HS65_LSS_XOR2X3 U17785 ( .A(n949), .B(n9682), .Z(n5955) );
  HS65_LSS_XNOR3X2 U17786 ( .A(n3216), .B(n5957), .C(n5958), .Z(n5956) );
  HS65_LSS_XOR3X2 U17787 ( .A(n2774), .B(n9200), .C(n2821), .Z(n5957) );
  HS65_LS_NOR2X2 U17788 ( .A(n9302), .B(n9319), .Z(n5751) );
  HS65_LS_NOR2X2 U17789 ( .A(n9381), .B(n9374), .Z(n7343) );
  HS65_LS_NOR2X2 U17790 ( .A(sa01[7]), .B(n9235), .Z(n7405) );
  HS65_LS_NOR2X2 U17791 ( .A(n9402), .B(n9236), .Z(n5813) );
  HS65_LS_NOR2X2 U17792 ( .A(n9385), .B(n9389), .Z(n5946) );
  HS65_LS_NOR2X2 U17793 ( .A(sa22[7]), .B(sa22[6]), .Z(n5887) );
  HS65_LS_NOR2X2 U17794 ( .A(n9390), .B(sa12[6]), .Z(n7538) );
  HS65_LS_NOR2X2 U17795 ( .A(n9305), .B(n9308), .Z(n7479) );
  HS65_LS_NOR2X2 U17796 ( .A(n602), .B(n9329), .Z(n9061) );
  HS65_LS_NOR2X2 U17797 ( .A(n115), .B(n9313), .Z(n9119) );
  HS65_LS_NOR2X2 U17798 ( .A(n44), .B(n9304), .Z(n5737) );
  HS65_LS_NOR2X2 U17799 ( .A(n570), .B(n9369), .Z(n7329) );
  HS65_LS_NOR2X2 U17800 ( .A(n490), .B(n9325), .Z(n5931) );
  HS65_LS_NOR2X2 U17801 ( .A(n271), .B(n9363), .Z(n5872) );
  HS65_LS_NOR2X2 U17802 ( .A(n708), .B(n9397), .Z(n5799) );
  HS65_LS_NOR2X2 U17803 ( .A(n178), .B(sa03[2]), .Z(n4156) );
  HS65_LS_NOR2X2 U17804 ( .A(n313), .B(n9303), .Z(n7523) );
  HS65_LS_NOR2X2 U17805 ( .A(n92), .B(sa23[2]), .Z(n7464) );
  HS65_LS_NOR2X2 U17806 ( .A(n526), .B(n9396), .Z(n7391) );
  HS65_LS_NOR2X2 U17807 ( .A(n229), .B(n9391), .Z(n4229) );
  HS65_LS_NOR2X2 U17808 ( .A(sa33[3]), .B(n9304), .Z(n5757) );
  HS65_LS_NOR2X2 U17809 ( .A(n9237), .B(n9369), .Z(n7349) );
  HS65_LS_NOR2X2 U17810 ( .A(n9354), .B(n9325), .Z(n5943) );
  HS65_LS_NOR2X2 U17811 ( .A(n9352), .B(n9363), .Z(n5884) );
  HS65_LS_NOR2X2 U17812 ( .A(n9321), .B(n9397), .Z(n5819) );
  HS65_LS_NOR2X2 U17813 ( .A(n9240), .B(n9303), .Z(n7535) );
  HS65_LS_NOR2X2 U17814 ( .A(sa23[3]), .B(sa23[2]), .Z(n7476) );
  HS65_LS_NOR2X2 U17815 ( .A(n9353), .B(n9396), .Z(n7411) );
  HS65_LS_NOR2X2 U17816 ( .A(n400), .B(n9376), .Z(n9002) );
  HS65_LS_NOR2X2 U17817 ( .A(n359), .B(n9243), .Z(n8934) );
  HS65_LS_NOR2X2 U17818 ( .A(sa20[1]), .B(n9384), .Z(n9038) );
  HS65_LS_NOR2X2 U17819 ( .A(n9241), .B(n9317), .Z(n9096) );
  HS65_LS_NOR2X2 U17820 ( .A(n340), .B(n9357), .Z(n8918) );
  HS65_LS_NOR2X2 U17821 ( .A(n385), .B(n9375), .Z(n8978) );
  HS65_LS_NOR2X2 U17822 ( .A(n427), .B(n9343), .Z(n4351) );
  HS65_LS_NOR2X2 U17823 ( .A(n207), .B(sa32[7]), .Z(n4230) );
  HS65_LS_NOR2X2 U17824 ( .A(n651), .B(n9383), .Z(n4287) );
  HS65_LS_NOR2AX3 U17825 ( .A(n9326), .B(n9346), .Z(n5945) );
  HS65_LS_NOR2AX3 U17826 ( .A(n9364), .B(n9362), .Z(n5886) );
  HS65_LS_NOR2AX3 U17827 ( .A(n9335), .B(n9345), .Z(n7537) );
  HS65_LS_NOR2AX3 U17828 ( .A(n9400), .B(n9320), .Z(n5824) );
  HS65_LS_NOR2AX3 U17829 ( .A(n9311), .B(n9306), .Z(n5762) );
  HS65_LS_NOR2AX3 U17830 ( .A(n9398), .B(sa23[4]), .Z(n7478) );
  HS65_LS_NOR2AX3 U17831 ( .A(n9367), .B(n9244), .Z(n7354) );
  HS65_LS_NOR2AX3 U17832 ( .A(n9395), .B(n9328), .Z(n7416) );
  HS65_LS_NOR2X2 U17833 ( .A(n9399), .B(n9347), .Z(n9044) );
  HS65_LS_NOR2X2 U17834 ( .A(n9309), .B(n9245), .Z(n9102) );
  HS65_LS_NOR2AX3 U17835 ( .A(n9330), .B(n9238), .Z(n4291) );
  HS65_LS_NOR2AX3 U17836 ( .A(n9316), .B(n9334), .Z(n4165) );
  HS65_LS_NOR2X2 U17837 ( .A(n9311), .B(n9306), .Z(n5750) );
  HS65_LS_NOR2X2 U17838 ( .A(n9367), .B(n9244), .Z(n7342) );
  HS65_LS_NOR2X2 U17839 ( .A(n9400), .B(n9320), .Z(n5812) );
  HS65_LS_NOR2X2 U17840 ( .A(n9326), .B(n9346), .Z(n5932) );
  HS65_LS_NOR2X2 U17841 ( .A(n9335), .B(n9345), .Z(n7524) );
  HS65_LS_NOR2X2 U17842 ( .A(n9398), .B(sa23[4]), .Z(n7465) );
  HS65_LS_NOR2X2 U17843 ( .A(n9395), .B(n9328), .Z(n7404) );
  HS65_LS_NOR2X2 U17844 ( .A(n9364), .B(n9362), .Z(n5873) );
  HS65_LS_IVX2 U17845 ( .A(n9394), .Z(n892) );
  HS65_LS_IVX2 U17846 ( .A(n9188), .Z(n810) );
  HS65_LS_IVX2 U17847 ( .A(n9174), .Z(n872) );
  HS65_LS_IVX2 U17848 ( .A(n9187), .Z(n911) );
  HS65_LS_IVX2 U17849 ( .A(n9173), .Z(n870) );
  HS65_LS_IVX2 U17850 ( .A(n9189), .Z(n829) );
  HS65_LS_IVX2 U17851 ( .A(n9191), .Z(n788) );
  HS65_LS_IVX2 U17852 ( .A(n9172), .Z(n891) );
  HS65_LS_IVX2 U17853 ( .A(n9393), .Z(n809) );
  HS65_LS_IVX2 U17854 ( .A(n9171), .Z(n811) );
  HS65_LS_IVX2 U17855 ( .A(n9386), .Z(n893) );
  HS65_LS_NOR2X2 U17856 ( .A(n911), .B(n9337), .Z(n2613) );
  HS65_LS_NOR2X2 U17857 ( .A(n829), .B(n9176), .Z(n1861) );
  HS65_LS_NOR2AX3 U17858 ( .A(n9326), .B(n470), .Z(n5934) );
  HS65_LS_NOR2AX3 U17859 ( .A(n9364), .B(n251), .Z(n5875) );
  HS65_LS_NOR2AX3 U17860 ( .A(n9335), .B(n293), .Z(n7526) );
  HS65_LS_NOR2AX3 U17861 ( .A(n9311), .B(n28), .Z(n5754) );
  HS65_LS_NOR2AX3 U17862 ( .A(n9398), .B(n72), .Z(n7467) );
  HS65_LS_NOR2AX3 U17863 ( .A(n9367), .B(n554), .Z(n7346) );
  HS65_LS_NOR2AX3 U17864 ( .A(n9400), .B(n692), .Z(n5816) );
  HS65_LS_NOR2AX3 U17865 ( .A(n9395), .B(n510), .Z(n7408) );
  HS65_LS_NOR2AX3 U17866 ( .A(n9316), .B(n184), .Z(n4155) );
  HS65_LS_NOR2AX3 U17867 ( .A(n9358), .B(n448), .Z(n4335) );
  HS65_LS_NOR2AX3 U17868 ( .A(n9376), .B(n400), .Z(n8994) );
  HS65_LS_NOR2AX3 U17869 ( .A(n9243), .B(n359), .Z(n8926) );
  HS65_LS_NOR2AX3 U17870 ( .A(n9307), .B(n50), .Z(n5738) );
  HS65_LS_NOR2AX3 U17871 ( .A(n9242), .B(n576), .Z(n7330) );
  HS65_LS_NOR2AX3 U17872 ( .A(n9349), .B(n492), .Z(n5921) );
  HS65_LS_NOR2AX3 U17873 ( .A(n9351), .B(n273), .Z(n5862) );
  HS65_LS_NOR2AX3 U17874 ( .A(n9239), .B(n315), .Z(n7513) );
  HS65_LS_NOR2AX3 U17875 ( .A(sa23[1]), .B(n94), .Z(n7454) );
  HS65_LS_NOR2AX3 U17876 ( .A(n9333), .B(n714), .Z(n5800) );
  HS65_LS_NOR2AX3 U17877 ( .A(n9332), .B(n532), .Z(n7392) );
  HS65_LS_IVX2 U17878 ( .A(n9182), .Z(n851) );
  HS65_LS_NOR2X2 U17879 ( .A(n9337), .B(n9187), .Z(n2618) );
  HS65_LS_NOR2X2 U17880 ( .A(n9167), .B(n9173), .Z(n1490) );
  HS65_LS_NOR2X2 U17881 ( .A(n9178), .B(n9191), .Z(n2242) );
  HS65_LS_NOR2X2 U17882 ( .A(n9176), .B(n9189), .Z(n1866) );
  HS65_LS_IVX2 U17883 ( .A(n9175), .Z(n890) );
  HS65_LS_IVX2 U17884 ( .A(n9186), .Z(n808) );
  HS65_LS_NOR2X2 U17885 ( .A(n790), .B(n9180), .Z(n2238) );
  HS65_LS_NOR2X2 U17886 ( .A(n831), .B(n9177), .Z(n1862) );
  HS65_LS_NOR2X2 U17887 ( .A(n913), .B(n9166), .Z(n2614) );
  HS65_LS_NOR2X2 U17888 ( .A(n872), .B(n9168), .Z(n1486) );
  HS65_LS_IVX2 U17889 ( .A(n9178), .Z(n789) );
  HS65_LS_IVX2 U17890 ( .A(n9168), .Z(n873) );
  HS65_LS_IVX2 U17891 ( .A(n9177), .Z(n832) );
  HS65_LS_IVX2 U17892 ( .A(n9167), .Z(n871) );
  HS65_LS_IVX2 U17893 ( .A(n9166), .Z(n914) );
  HS65_LS_IVX2 U17894 ( .A(n9180), .Z(n791) );
  HS65_LS_NOR2X2 U17895 ( .A(n871), .B(n9173), .Z(n1467) );
  HS65_LS_NOR2X2 U17896 ( .A(n912), .B(n9187), .Z(n2595) );
  HS65_LS_NOR2X2 U17897 ( .A(n789), .B(n9191), .Z(n2219) );
  HS65_LS_NOR2X2 U17898 ( .A(n830), .B(n9189), .Z(n1843) );
  HS65_LS_NOR2X2 U17899 ( .A(n870), .B(n9167), .Z(n1485) );
  HS65_LS_NOR2X2 U17900 ( .A(n788), .B(n9178), .Z(n2237) );
  HS65_LS_IVX2 U17901 ( .A(n9170), .Z(n933) );
  HS65_LS_IVX2 U17902 ( .A(n9169), .Z(n913) );
  HS65_LS_IVX2 U17903 ( .A(n9184), .Z(n831) );
  HS65_LS_IVX2 U17904 ( .A(n9339), .Z(n850) );
  HS65_LS_IVX2 U17905 ( .A(n9181), .Z(n932) );
  HS65_LS_IVX2 U17906 ( .A(n9338), .Z(n852) );
  HS65_LS_IVX2 U17907 ( .A(n9176), .Z(n830) );
  HS65_LS_IVX2 U17908 ( .A(n9337), .Z(n912) );
  HS65_LS_IVX2 U17909 ( .A(n9183), .Z(n934) );
  HS65_LS_IVX2 U17910 ( .A(n9185), .Z(n849) );
  HS65_LS_IVX2 U17911 ( .A(n9179), .Z(n931) );
  HS65_LS_NOR2X2 U17912 ( .A(sa32[7]), .B(n9368), .Z(n4227) );
  HS65_LS_NOR2X2 U17913 ( .A(n183), .B(sa03[3]), .Z(n4157) );
  HS65_LS_NOR2AX3 U17914 ( .A(sa20[1]), .B(n9384), .Z(n9055) );
  HS65_LS_NOR2AX3 U17915 ( .A(n9241), .B(n9317), .Z(n9113) );
  HS65_LS_NOR2AX3 U17916 ( .A(n9307), .B(n9300), .Z(n5760) );
  HS65_LS_NOR2AX3 U17917 ( .A(n9242), .B(n9372), .Z(n7352) );
  HS65_LS_NOR2X2 U17918 ( .A(n492), .B(n9349), .Z(n5939) );
  HS65_LS_NOR2X2 U17919 ( .A(n273), .B(n9351), .Z(n5880) );
  HS65_LS_NOR2X2 U17920 ( .A(n315), .B(n9239), .Z(n7531) );
  HS65_LS_NOR2X2 U17921 ( .A(n94), .B(sa23[1]), .Z(n7472) );
  HS65_LS_NOR2X2 U17922 ( .A(n714), .B(n9333), .Z(n5818) );
  HS65_LS_NOR2X2 U17923 ( .A(n532), .B(n9332), .Z(n7410) );
  HS65_LS_NOR2X2 U17924 ( .A(n9342), .B(n9322), .Z(n9037) );
  HS65_LS_NOR2X2 U17925 ( .A(n9247), .B(sa13[2]), .Z(n9095) );
  HS65_LS_NOR2X2 U17926 ( .A(sa32[1]), .B(n9391), .Z(n4219) );
  HS65_LS_NOR2X2 U17927 ( .A(n9350), .B(n9378), .Z(n4353) );
  HS65_LS_NOR2X2 U17928 ( .A(n9334), .B(n9316), .Z(n4158) );
  HS65_LS_NOR2X2 U17929 ( .A(n9238), .B(n9330), .Z(n4294) );
  HS65_LS_NOR2X2 U17930 ( .A(n184), .B(n9316), .Z(n4167) );
  HS65_LS_NOR2X2 U17931 ( .A(n9349), .B(n9380), .Z(n5941) );
  HS65_LS_NOR2X2 U17932 ( .A(n9351), .B(n9379), .Z(n5882) );
  HS65_LS_NOR2X2 U17933 ( .A(n9333), .B(n9312), .Z(n5815) );
  HS65_LS_NOR2X2 U17934 ( .A(n9239), .B(n9318), .Z(n7533) );
  HS65_LS_NOR2X2 U17935 ( .A(sa23[1]), .B(n9301), .Z(n7474) );
  HS65_LS_NOR2X2 U17936 ( .A(n9332), .B(n9392), .Z(n7407) );
  HS65_LS_NOR2X2 U17937 ( .A(n673), .B(n9327), .Z(n4292) );
  HS65_LS_NOR2X2 U17938 ( .A(n626), .B(n9342), .Z(n9050) );
  HS65_LS_NOR2X2 U17939 ( .A(n139), .B(n9247), .Z(n9108) );
  HS65_LS_NOR2AX3 U17940 ( .A(n9377), .B(n9361), .Z(n4220) );
  HS65_LS_NOR2AX3 U17941 ( .A(n9358), .B(n9341), .Z(n4349) );
  HS65_LS_NOR2X2 U17942 ( .A(n9299), .B(n9298), .Z(n4160) );
  HS65_LS_NOR2X2 U17943 ( .A(n360), .B(n9370), .Z(n8927) );
  HS65_LS_NOR2X2 U17944 ( .A(n406), .B(n9360), .Z(n9001) );
  HS65_LS_NOR2X2 U17945 ( .A(n209), .B(n9387), .Z(n4211) );
  HS65_LS_NOR2X2 U17946 ( .A(n627), .B(sa20[1]), .Z(n9051) );
  HS65_LS_NOR2X2 U17947 ( .A(n140), .B(n9241), .Z(n9109) );
  HS65_LS_NOR2X2 U17948 ( .A(n450), .B(n9350), .Z(n4348) );
  HS65_LS_NOR2X2 U17949 ( .A(n230), .B(sa32[1]), .Z(n4224) );
  HS65_LSS_XNOR2X3 U17950 ( .A(n2510), .B(n9225), .Z(n1016) );
  HS65_LS_NOR4ABX2 U17951 ( .A(n2511), .B(n2512), .C(n2513), .D(n2514), .Z(
        n2510) );
  HS65_LS_CBI4I1X3 U17952 ( .A(n2329), .B(n2257), .C(n2283), .D(n2462), .Z(
        n2514) );
  HS65_LS_CBI4I6X2 U17953 ( .A(n901), .B(n2484), .C(n922), .D(n2533), .Z(n2511) );
  HS65_LSS_XNOR2X3 U17954 ( .A(n1913), .B(n9215), .Z(n1005) );
  HS65_LS_NOR3X1 U17955 ( .A(n1914), .B(n1915), .C(n1916), .Z(n1913) );
  HS65_LS_NAND4ABX3 U17956 ( .A(n1941), .B(n1942), .C(n1943), .D(n1944), .Z(
        n1914) );
  HS65_LS_OAI212X3 U17957 ( .A(n1881), .B(n1886), .C(n1908), .D(n1938), .E(
        n1939), .Z(n1915) );
  HS65_LSS_XOR2X3 U17958 ( .A(n1016), .B(n9213), .Z(n1112) );
  HS65_LSS_XOR2X3 U17959 ( .A(n1013), .B(n9212), .Z(n1109) );
  HS65_LSS_XNOR2X3 U17960 ( .A(n1954), .B(n9214), .Z(n1006) );
  HS65_LS_NOR3X1 U17961 ( .A(n1955), .B(n1956), .C(n1957), .Z(n1954) );
  HS65_LS_OAI212X3 U17962 ( .A(n1958), .B(n1882), .C(n1959), .D(n1960), .E(
        n1961), .Z(n1957) );
  HS65_LS_NAND4ABX3 U17963 ( .A(n1962), .B(n1963), .C(n1964), .D(n1965), .Z(
        n1956) );
  HS65_LSS_XNOR2X3 U17964 ( .A(n1578), .B(n9211), .Z(n998) );
  HS65_LS_NOR3X1 U17965 ( .A(n1579), .B(n1580), .C(n1581), .Z(n1578) );
  HS65_LS_OAI212X3 U17966 ( .A(n1582), .B(n1506), .C(n1583), .D(n1584), .E(
        n1585), .Z(n1581) );
  HS65_LS_NAND4ABX3 U17967 ( .A(n1586), .B(n1587), .C(n1588), .D(n1589), .Z(
        n1580) );
  HS65_LSS_XOR2X3 U17968 ( .A(n1008), .B(n9210), .Z(n1104) );
  HS65_LSS_XOR2X3 U17969 ( .A(n1005), .B(n9209), .Z(n1101) );
  HS65_LSS_XOR2X3 U17970 ( .A(n1006), .B(n9208), .Z(n1102) );
  HS65_LSS_XOR2X3 U17971 ( .A(n1014), .B(n9207), .Z(n1110) );
  HS65_LSS_XOR2X3 U17972 ( .A(n998), .B(n9206), .Z(n1094) );
  HS65_LSS_XNOR2X3 U17973 ( .A(n9282), .B(n1114), .Z(n1082) );
  HS65_LSS_XNOR2X3 U17974 ( .A(n9280), .B(n1091), .Z(n1036) );
  HS65_LSS_XNOR2X3 U17975 ( .A(n9287), .B(n1109), .Z(n1072) );
  HS65_LSS_XNOR2X3 U17976 ( .A(n9250), .B(n1092), .Z(n1038) );
  HS65_LS_NOR2AX3 U17977 ( .A(n9377), .B(n224), .Z(n4226) );
  HS65_LSS_XNOR2X3 U17978 ( .A(n9271), .B(n1518), .Z(n996) );
  HS65_LS_NAND4ABX3 U17979 ( .A(n1519), .B(n1520), .C(n1521), .D(n1522), .Z(
        n1518) );
  HS65_LS_CBI4I1X3 U17980 ( .A(n1534), .B(n1504), .C(n1535), .D(n1536), .Z(
        n1519) );
  HS65_LS_CBI4I1X3 U17981 ( .A(n1530), .B(n1531), .C(n1532), .D(n1533), .Z(
        n1520) );
  HS65_LSS_XNOR2X3 U17982 ( .A(n9297), .B(n1106), .Z(n1066) );
  HS65_LSS_XNOR2X3 U17983 ( .A(n9292), .B(n1112), .Z(n1078) );
  HS65_LSS_XNOR2X3 U17984 ( .A(n9281), .B(n1090), .Z(n1034) );
  HS65_LSS_XNOR2X3 U17985 ( .A(n9291), .B(n1108), .Z(n1070) );
  HS65_LSS_XNOR2X3 U17986 ( .A(n9258), .B(n2183), .Z(n1010) );
  HS65_LS_NAND4ABX3 U17987 ( .A(n2184), .B(n2185), .C(n2186), .D(n2187), .Z(
        n2183) );
  HS65_LS_MX41X4 U17988 ( .D0(n784), .S0(n801), .D1(n785), .S1(n793), .D2(n804), .S2(n777), .D3(n805), .S3(n1930), .Z(n2185) );
  HS65_LS_NOR4ABX2 U17989 ( .A(n1928), .B(n2063), .C(n2188), .D(n2077), .Z(
        n2187) );
  HS65_LSS_XNOR2X3 U17990 ( .A(n9263), .B(n2243), .Z(n1011) );
  HS65_LS_NAND4ABX3 U17991 ( .A(n2244), .B(n2245), .C(n2246), .D(n2247), .Z(
        n2243) );
  HS65_LS_OAI212X3 U17992 ( .A(n2255), .B(n2256), .C(n2257), .D(n2258), .E(
        n2259), .Z(n2245) );
  HS65_LS_NAND4ABX3 U17993 ( .A(n2265), .B(n2266), .C(n2267), .D(n2268), .Z(
        n2244) );
  HS65_LSS_XNOR2X3 U17994 ( .A(n9257), .B(n2559), .Z(n1018) );
  HS65_LS_NAND4ABX3 U17995 ( .A(n2560), .B(n2561), .C(n2562), .D(n2563), .Z(
        n2559) );
  HS65_LS_NOR4ABX2 U17996 ( .A(n2304), .B(n2439), .C(n2564), .D(n2453), .Z(
        n2563) );
  HS65_LS_MX41X4 U17997 ( .D0(n907), .S0(n924), .D1(n908), .S1(n916), .D2(n927), .S2(n900), .D3(n928), .S3(n2306), .Z(n2561) );
  HS65_LSS_XNOR2X3 U17998 ( .A(n9268), .B(n2270), .Z(n1012) );
  HS65_LS_NAND4ABX3 U17999 ( .A(n2271), .B(n2272), .C(n2273), .D(n2274), .Z(
        n2270) );
  HS65_LS_CBI4I1X3 U18000 ( .A(n2286), .B(n2256), .C(n2287), .D(n2288), .Z(
        n2271) );
  HS65_LS_CBI4I1X3 U18001 ( .A(n2282), .B(n2283), .C(n2284), .D(n2285), .Z(
        n2272) );
  HS65_LSS_XNOR2X3 U18002 ( .A(n9289), .B(n1110), .Z(n1074) );
  HS65_LSS_XNOR2X3 U18003 ( .A(n9283), .B(n1083), .Z(n1020) );
  HS65_LSS_XNOR2X3 U18004 ( .A(n9295), .B(n1104), .Z(n1062) );
  HS65_LSS_XNOR2X3 U18005 ( .A(n9288), .B(n1102), .Z(n1058) );
  HS65_LSS_XNOR2X3 U18006 ( .A(n9286), .B(n1101), .Z(n1056) );
  HS65_LSS_XNOR2X3 U18007 ( .A(n9296), .B(n1111), .Z(n1076) );
  HS65_LSS_XNOR2X3 U18008 ( .A(n9275), .B(n1085), .Z(n1024) );
  HS65_LSS_XNOR2X3 U18009 ( .A(n9284), .B(n1100), .Z(n1054) );
  HS65_LSS_XNOR2X3 U18010 ( .A(n9276), .B(n1086), .Z(n1026) );
  HS65_LSS_XNOR2X3 U18011 ( .A(n9293), .B(n1105), .Z(n1064) );
  HS65_LSS_XNOR2X3 U18012 ( .A(n9290), .B(n1103), .Z(n1060) );
  HS65_LSS_XNOR2X3 U18013 ( .A(n9285), .B(n1113), .Z(n1080) );
  HS65_LSS_XNOR2X3 U18014 ( .A(n9254), .B(n1099), .Z(n1052) );
  HS65_LSS_XNOR2X3 U18015 ( .A(n9279), .B(n1089), .Z(n1032) );
  HS65_LSS_XNOR2X3 U18016 ( .A(n9251), .B(n1094), .Z(n1042) );
  HS65_LSS_XNOR2X3 U18017 ( .A(n9264), .B(n2158), .Z(n1009) );
  HS65_LS_NAND4ABX3 U18018 ( .A(n2159), .B(n2160), .C(n2161), .D(n2162), .Z(
        n2158) );
  HS65_LS_AOI222X2 U18019 ( .A(n795), .B(n773), .C(n792), .D(n2181), .E(n804), 
        .F(n772), .Z(n2161) );
  HS65_LS_CB4I6X4 U18020 ( .A(n776), .B(n781), .C(n803), .D(n2079), .Z(n2159)
         );
  HS65_LSS_XNOR2X3 U18021 ( .A(n9269), .B(n2017), .Z(n1007) );
  HS65_LS_NAND4ABX3 U18022 ( .A(n2018), .B(n2019), .C(n2020), .D(n2021), .Z(
        n2017) );
  HS65_LS_MX41X4 U18023 ( .D0(n774), .S0(n798), .D1(n802), .S1(n786), .D2(n772), .S2(n793), .D3(n804), .S3(n1930), .Z(n2019) );
  HS65_LS_AOI212X2 U18024 ( .A(n787), .B(n2022), .C(n803), .D(n1999), .E(n2023), .Z(n2021) );
  HS65_LSS_XNOR2X3 U18025 ( .A(n9234), .B(n994), .Z(n1090) );
  HS65_LSS_XNOR2X3 U18026 ( .A(n9233), .B(n996), .Z(n1092) );
  HS65_LSS_XNOR2X3 U18027 ( .A(n9230), .B(n1002), .Z(n1098) );
  HS65_LSS_XNOR2X3 U18028 ( .A(n9229), .B(n1011), .Z(n1107) );
  HS65_LSS_XNOR2X3 U18029 ( .A(n9232), .B(n1010), .Z(n1106) );
  HS65_LSS_XNOR2X3 U18030 ( .A(n9231), .B(n995), .Z(n1091) );
  HS65_LSS_XNOR2X3 U18031 ( .A(n9228), .B(n1018), .Z(n1114) );
  HS65_LSS_XNOR2X3 U18032 ( .A(n9227), .B(n1012), .Z(n1108) );
  HS65_LSS_XNOR2X3 U18033 ( .A(n9220), .B(n991), .Z(n1087) );
  HS65_LSS_XNOR2X3 U18034 ( .A(n9219), .B(n1001), .Z(n1097) );
  HS65_LSS_XNOR2X3 U18035 ( .A(n9218), .B(n999), .Z(n1095) );
  HS65_LSS_XNOR2X3 U18036 ( .A(n9224), .B(n1004), .Z(n1100) );
  HS65_LSS_XNOR2X3 U18037 ( .A(n9223), .B(n1017), .Z(n1113) );
  HS65_LSS_XNOR2X3 U18038 ( .A(n9222), .B(n1015), .Z(n1111) );
  HS65_LSS_XNOR2X3 U18039 ( .A(n9221), .B(n1009), .Z(n1105) );
  HS65_LS_NOR2X2 U18040 ( .A(n50), .B(n9307), .Z(n5756) );
  HS65_LS_NOR2X2 U18041 ( .A(n576), .B(n9242), .Z(n7348) );
  HS65_LSS_XNOR2X3 U18042 ( .A(n9217), .B(n1003), .Z(n1099) );
  HS65_LSS_XNOR2X3 U18043 ( .A(n9216), .B(n1007), .Z(n1103) );
  HS65_LS_NOR2X2 U18044 ( .A(n161), .B(n9298), .Z(n4161) );
  HS65_LS_NOR2X2 U18045 ( .A(n27), .B(n9302), .Z(n5755) );
  HS65_LS_NOR2X2 U18046 ( .A(n553), .B(n9381), .Z(n7347) );
  HS65_LS_NOR2X2 U18047 ( .A(n71), .B(n9305), .Z(n7477) );
  HS65_LS_NOR2X2 U18048 ( .A(n469), .B(n9385), .Z(n5944) );
  HS65_LS_NOR2X2 U18049 ( .A(n292), .B(n9390), .Z(n7536) );
  HS65_LS_NOR2X2 U18050 ( .A(n250), .B(sa22[7]), .Z(n5885) );
  HS65_LS_NOR2X2 U18051 ( .A(n691), .B(n9402), .Z(n5817) );
  HS65_LS_NOR2X2 U18052 ( .A(n509), .B(sa01[7]), .Z(n7409) );
  HS65_LS_NOR2X2 U18053 ( .A(n575), .B(n9237), .Z(n7344) );
  HS65_LS_NOR2X2 U18054 ( .A(n49), .B(sa33[3]), .Z(n5752) );
  HS65_LS_NOR2X2 U18055 ( .A(n491), .B(n9354), .Z(n5920) );
  HS65_LS_NOR2X2 U18056 ( .A(n272), .B(n9352), .Z(n5861) );
  HS65_LS_NOR2X2 U18057 ( .A(n314), .B(n9240), .Z(n7512) );
  HS65_LS_NOR2X2 U18058 ( .A(n93), .B(sa23[3]), .Z(n7453) );
  HS65_LS_NOR2X2 U18059 ( .A(n713), .B(n9321), .Z(n5814) );
  HS65_LS_NOR2X2 U18060 ( .A(n531), .B(n9353), .Z(n7406) );
  HS65_LSS_XNOR2X3 U18061 ( .A(n9205), .B(n987), .Z(n1083) );
  HS65_LSS_XNOR2X3 U18062 ( .A(n9204), .B(n993), .Z(n1089) );
  HS65_LSS_XNOR2X3 U18063 ( .A(n9203), .B(n988), .Z(n1084) );
  HS65_LSS_XOR2X3 U18064 ( .A(n2330), .B(n954), .Z(n1014) );
  HS65_LS_NOR3X1 U18065 ( .A(n2331), .B(n2332), .C(n2333), .Z(n2330) );
  HS65_LS_OAI212X3 U18066 ( .A(n2334), .B(n2258), .C(n2335), .D(n2336), .E(
        n2337), .Z(n2333) );
  HS65_LS_NAND4ABX3 U18067 ( .A(n2338), .B(n2339), .C(n2340), .D(n2341), .Z(
        n2332) );
  HS65_LSS_XOR2X3 U18068 ( .A(n3016), .B(n9234), .Z(n9757) );
  HS65_LSS_XNOR2X3 U18069 ( .A(n2816), .B(n9280), .Z(n9790) );
  HS65_LSS_XNOR2X3 U18070 ( .A(n2815), .B(n9250), .Z(n9791) );
  HS65_LSS_XNOR2X3 U18071 ( .A(n2823), .B(n9233), .Z(n9759) );
  HS65_LSS_XNOR2X3 U18072 ( .A(n2831), .B(n9271), .Z(n9727) );
  HS65_LSS_XNOR2X3 U18073 ( .A(n2766), .B(n9287), .Z(n9808) );
  HS65_LSS_XNOR2X3 U18074 ( .A(n2761), .B(n9282), .Z(n9813) );
  HS65_LSS_XOR2X3 U18075 ( .A(n2832), .B(n9261), .Z(n9726) );
  HS65_LSS_XOR2X3 U18076 ( .A(n2763), .B(n9292), .Z(n9811) );
  HS65_LSS_XOR2X3 U18077 ( .A(n2785), .B(n9297), .Z(n9805) );
  HS65_LSS_XOR2X3 U18078 ( .A(n2824), .B(n9231), .Z(n9758) );
  HS65_LSS_XOR2X3 U18079 ( .A(n2801), .B(n9258), .Z(n9741) );
  HS65_LSS_XOR2X3 U18080 ( .A(n2793), .B(n9232), .Z(n9773) );
  HS65_LSS_XOR2X3 U18081 ( .A(n2817), .B(n9230), .Z(n9765) );
  HS65_LSS_XOR2X3 U18082 ( .A(n2776), .B(n9229), .Z(n9774) );
  HS65_LSS_XOR2X3 U18083 ( .A(n2784), .B(n9263), .Z(n9742) );
  HS65_LSS_XNOR2X3 U18084 ( .A(n2775), .B(n9227), .Z(n9775) );
  HS65_LSS_XNOR2X3 U18085 ( .A(n2783), .B(n9268), .Z(n9743) );
  HS65_LSS_XNOR2X3 U18086 ( .A(n2769), .B(n9228), .Z(n9781) );
  HS65_LSS_XNOR2X3 U18087 ( .A(n2777), .B(n9257), .Z(n9749) );
  HS65_LSS_XOR2X3 U18088 ( .A(n2774), .B(n9212), .Z(n9776) );
  HS65_LSS_XOR2X3 U18089 ( .A(n2771), .B(n9213), .Z(n9779) );
  HS65_LSS_XNOR2X3 U18090 ( .A(n2767), .B(n9291), .Z(n9807) );
  HS65_LSS_XOR2X3 U18091 ( .A(n2782), .B(n9226), .Z(n9744) );
  HS65_LSS_XOR2X3 U18092 ( .A(n2908), .B(n9281), .Z(n9789) );
  HS65_LSS_XOR2X3 U18093 ( .A(n2779), .B(n9225), .Z(n9747) );
  HS65_LSS_XOR2X3 U18094 ( .A(n3015), .B(n9283), .Z(n9782) );
  HS65_LSS_XOR2X3 U18095 ( .A(n2799), .B(n9224), .Z(n9767) );
  HS65_LSS_XOR2X3 U18096 ( .A(n2787), .B(n9295), .Z(n9803) );
  HS65_LSS_XNOR2X3 U18097 ( .A(n2791), .B(n9284), .Z(n9799) );
  HS65_LSS_XNOR2X3 U18098 ( .A(n3013), .B(n9275), .Z(n9784) );
  HS65_LSS_XOR2X3 U18099 ( .A(n2764), .B(n9296), .Z(n9810) );
  HS65_LSS_XOR2X3 U18100 ( .A(n2770), .B(n9223), .Z(n9780) );
  HS65_LSS_XOR2X3 U18101 ( .A(n2798), .B(n9209), .Z(n9768) );
  HS65_LSS_XOR2X3 U18102 ( .A(n2795), .B(n9210), .Z(n9771) );
  HS65_LSS_XNOR2X3 U18103 ( .A(n2772), .B(n9222), .Z(n9778) );
  HS65_LSS_XNOR2X3 U18104 ( .A(n2797), .B(n9208), .Z(n9769) );
  HS65_LSS_XOR2X3 U18105 ( .A(n2806), .B(n9215), .Z(n9736) );
  HS65_LSS_XNOR2X3 U18106 ( .A(n2773), .B(n9207), .Z(n9777) );
  HS65_LSS_XOR2X3 U18107 ( .A(n3019), .B(n9220), .Z(n9754) );
  HS65_LSS_XOR2X3 U18108 ( .A(n2818), .B(n9219), .Z(n9764) );
  HS65_LSS_XOR2X3 U18109 ( .A(n2820), .B(n9218), .Z(n9762) );
  HS65_LSS_XOR2X3 U18110 ( .A(n2786), .B(n9293), .Z(n9804) );
  HS65_LSS_XOR2X3 U18111 ( .A(n2794), .B(n9221), .Z(n9772) );
  HS65_LSS_XOR2X3 U18112 ( .A(n2802), .B(n9264), .Z(n9740) );
  HS65_LSS_XOR2X3 U18113 ( .A(n2788), .B(n9290), .Z(n9802) );
  HS65_LSS_XOR2X3 U18114 ( .A(n2762), .B(n9285), .Z(n9812) );
  HS65_LSS_XOR2X3 U18115 ( .A(n2669), .B(n9169), .Z(n9819) );
  HS65_LSS_XOR2X3 U18116 ( .A(n2640), .B(n9170), .Z(n9815) );
  HS65_LSS_XOR2X3 U18117 ( .A(n2717), .B(n9184), .Z(n9835) );
  HS65_LSS_XNOR2X3 U18118 ( .A(n2805), .B(n9214), .Z(n9737) );
  HS65_LSS_XNOR2X3 U18119 ( .A(n2813), .B(n9251), .Z(n9793) );
  HS65_LSS_XNOR2X3 U18120 ( .A(n2630), .B(n9279), .Z(n9788) );
  HS65_LSS_XNOR2X3 U18121 ( .A(n2796), .B(n9216), .Z(n9770) );
  HS65_LSS_XNOR2X3 U18122 ( .A(n2804), .B(n9269), .Z(n9738) );
  HS65_LSS_XOR2X3 U18123 ( .A(n2821), .B(n9206), .Z(n9761) );
  HS65_LSS_XOR2X3 U18124 ( .A(n2792), .B(n9254), .Z(n9798) );
  HS65_LSS_XOR2X3 U18125 ( .A(n2800), .B(n9217), .Z(n9766) );
  HS65_LSS_XOR2X3 U18126 ( .A(n2829), .B(n9211), .Z(n9729) );
  HS65_LSS_XOR2X3 U18127 ( .A(n2653), .B(n9179), .Z(n9817) );
  HS65_LSS_XOR2X3 U18128 ( .A(n2707), .B(n9185), .Z(n9833) );
  HS65_LSS_XOR2X3 U18129 ( .A(n2691), .B(n9183), .Z(n9814) );
  HS65_LSS_XOR2X3 U18130 ( .A(n2701), .B(n9339), .Z(n9832) );
  HS65_LSS_XOR2X3 U18131 ( .A(n2646), .B(n9181), .Z(n9816) );
  HS65_LSS_XOR2X3 U18132 ( .A(n2722), .B(n9176), .Z(n9836) );
  HS65_LSS_XOR2X3 U18133 ( .A(n2907), .B(n9337), .Z(n9820) );
  HS65_LSS_XOR2X3 U18134 ( .A(n2728), .B(n9338), .Z(n9830) );
  HS65_LSS_XNOR2X3 U18135 ( .A(n2289), .B(n9226), .Z(n1013) );
  HS65_LS_NOR3X1 U18136 ( .A(n2290), .B(n2291), .C(n2292), .Z(n2289) );
  HS65_LS_NAND4ABX3 U18137 ( .A(n2317), .B(n2318), .C(n2319), .D(n2320), .Z(
        n2290) );
  HS65_LS_OAI212X3 U18138 ( .A(n2257), .B(n2262), .C(n2284), .D(n2314), .E(
        n2315), .Z(n2291) );
  HS65_LSS_XOR2X3 U18139 ( .A(n3017), .B(n9204), .Z(n9756) );
  HS65_LSS_XOR2X3 U18140 ( .A(n3219), .B(n9205), .Z(n9750) );
  HS65_LSS_XNOR2X3 U18141 ( .A(n9276), .B(n3012), .Z(n9785) );
  HS65_LSS_XOR2X3 U18142 ( .A(n2680), .B(n9173), .Z(n9829) );
  HS65_LSS_XOR2X3 U18143 ( .A(n2667), .B(n9174), .Z(n9827) );
  HS65_LSS_XOR2X3 U18144 ( .A(n2645), .B(n9188), .Z(n9839) );
  HS65_LSS_XOR2X3 U18145 ( .A(n2736), .B(n9394), .Z(n9823) );
  HS65_LSS_XOR2X3 U18146 ( .A(n2687), .B(n9191), .Z(n9845) );
  HS65_LSS_XOR2X3 U18147 ( .A(n2682), .B(n9187), .Z(n9821) );
  HS65_LSS_XOR2X3 U18148 ( .A(n2696), .B(n9182), .Z(n9831) );
  HS65_LSS_XOR2X3 U18149 ( .A(n2727), .B(n9189), .Z(n9837) );
  HS65_LSS_XOR2X3 U18150 ( .A(n2757), .B(n9167), .Z(n9828) );
  HS65_LSS_XOR2X3 U18151 ( .A(n2660), .B(n9168), .Z(n9826) );
  HS65_LSS_XOR2X3 U18152 ( .A(n2681), .B(n9178), .Z(n9844) );
  HS65_LSS_XOR2X3 U18153 ( .A(n2659), .B(n9166), .Z(n9818) );
  HS65_LSS_XOR2X3 U18154 ( .A(n2639), .B(n9386), .Z(n9822) );
  HS65_LSS_XOR2X3 U18155 ( .A(n2668), .B(n9180), .Z(n9842) );
  HS65_LSS_XOR2X3 U18156 ( .A(n2712), .B(n9177), .Z(n9834) );
  HS65_LSS_XOR2X3 U18157 ( .A(n2732), .B(n9171), .Z(n9838) );
  HS65_LSS_XOR2X3 U18158 ( .A(n3220), .B(n9260), .Z(n9725) );
  HS65_LSS_XOR2X3 U18159 ( .A(n3218), .B(n9203), .Z(n9751) );
  HS65_LSS_XOR2X3 U18160 ( .A(n2827), .B(n9195), .Z(n9731) );
  HS65_LSS_XOR2X3 U18161 ( .A(n2819), .B(n9201), .Z(n9763) );
  HS65_LSS_XOR2X3 U18162 ( .A(n2811), .B(n9255), .Z(n9795) );
  HS65_LS_IVX2 U18163 ( .A(sa02[6]), .Z(n338) );
  HS65_LS_IVX2 U18164 ( .A(n9310), .Z(n164) );
  HS65_LS_IVX2 U18165 ( .A(n9365), .Z(n427) );
  HS65_LS_IVX2 U18166 ( .A(n9356), .Z(n340) );
  HS65_LS_IVX2 U18167 ( .A(n9370), .Z(n361) );
  HS65_LS_IVX2 U18168 ( .A(n9347), .Z(n605) );
  HS65_LS_IVX2 U18169 ( .A(n9373), .Z(n383) );
  HS65_LS_IVX2 U18170 ( .A(n9245), .Z(n118) );
  HS65_LS_IVX2 U18171 ( .A(sa13[2]), .Z(n139) );
  HS65_LS_IVX2 U18172 ( .A(n9322), .Z(n626) );
  HS65_LS_IVX2 U18173 ( .A(n9388), .Z(n651) );
  HS65_LS_IVX2 U18174 ( .A(n9325), .Z(n491) );
  HS65_LS_IVX2 U18175 ( .A(n9363), .Z(n272) );
  HS65_LS_IVX2 U18176 ( .A(n9304), .Z(n49) );
  HS65_LS_IVX2 U18177 ( .A(n9378), .Z(n450) );
  HS65_LS_IVX2 U18178 ( .A(n9324), .Z(n673) );
  HS65_LS_IVX2 U18179 ( .A(n9391), .Z(n230) );
  HS65_LS_IVX2 U18180 ( .A(n9368), .Z(n207) );
  HS65_LS_IVX2 U18181 ( .A(n9298), .Z(n162) );
  HS65_LS_IVX2 U18182 ( .A(n9348), .Z(n385) );
  HS65_LS_IVX2 U18183 ( .A(n9303), .Z(n314) );
  HS65_LS_IVX2 U18184 ( .A(sa23[2]), .Z(n93) );
  HS65_LS_IVX2 U18185 ( .A(n9369), .Z(n575) );
  HS65_LS_IVX2 U18186 ( .A(n9371), .Z(n406) );
  HS65_LS_IVX2 U18187 ( .A(n9397), .Z(n713) );
  HS65_LS_IVX2 U18188 ( .A(n9396), .Z(n531) );
  HS65_LS_IVX2 U18189 ( .A(n9387), .Z(n208) );
  HS65_LS_IVX2 U18190 ( .A(n9359), .Z(n428) );
  HS65_LS_IVX2 U18191 ( .A(n9323), .Z(n652) );
  HS65_LS_IVX2 U18192 ( .A(sa03[3]), .Z(n178) );
  HS65_LS_IVX2 U18193 ( .A(n9246), .Z(n602) );
  HS65_LS_IVX2 U18194 ( .A(n9314), .Z(n115) );
  HS65_LS_IVX2 U18195 ( .A(n9306), .Z(n28) );
  HS65_LS_IVX2 U18196 ( .A(n9384), .Z(n627) );
  HS65_LS_IVX2 U18197 ( .A(n9244), .Z(n554) );
  HS65_LS_IVX2 U18198 ( .A(n9346), .Z(n470) );
  HS65_LS_IVX2 U18199 ( .A(n9389), .Z(n469) );
  HS65_LS_IVX2 U18200 ( .A(n9380), .Z(n492) );
  HS65_LS_IVX2 U18201 ( .A(n9362), .Z(n251) );
  HS65_LS_IVX2 U18202 ( .A(sa22[6]), .Z(n250) );
  HS65_LS_IVX2 U18203 ( .A(n9379), .Z(n273) );
  HS65_LS_IVX2 U18204 ( .A(n9320), .Z(n692) );
  HS65_LS_IVX2 U18205 ( .A(n9300), .Z(n50) );
  HS65_LS_IVX2 U18206 ( .A(n9319), .Z(n27) );
  HS65_LS_IVX2 U18207 ( .A(n9317), .Z(n140) );
  HS65_LS_IVX2 U18208 ( .A(n9345), .Z(n293) );
  HS65_LS_IVX2 U18209 ( .A(sa12[6]), .Z(n292) );
  HS65_LS_IVX2 U18210 ( .A(n9318), .Z(n315) );
  HS65_LS_IVX2 U18211 ( .A(sa23[4]), .Z(n72) );
  HS65_LS_IVX2 U18212 ( .A(n9301), .Z(n94) );
  HS65_LS_IVX2 U18213 ( .A(n9308), .Z(n71) );
  HS65_LS_IVX2 U18214 ( .A(n9372), .Z(n576) );
  HS65_LS_IVX2 U18215 ( .A(n9374), .Z(n553) );
  HS65_LS_IVX2 U18216 ( .A(n9328), .Z(n510) );
  HS65_LS_IVX2 U18217 ( .A(n9312), .Z(n714) );
  HS65_LS_IVX2 U18218 ( .A(n9235), .Z(n509) );
  HS65_LS_IVX2 U18219 ( .A(n9236), .Z(n691) );
  HS65_LS_IVX2 U18220 ( .A(n9392), .Z(n532) );
  HS65_LS_IVX2 U18221 ( .A(n9341), .Z(n448) );
  HS65_LS_IVX2 U18222 ( .A(n9238), .Z(n674) );
  HS65_LS_IVX2 U18223 ( .A(n9361), .Z(n224) );
  HS65_LS_IVX2 U18224 ( .A(n9401), .Z(n400) );
  HS65_LS_IVX2 U18225 ( .A(n9336), .Z(n359) );
  HS65_LS_IVX2 U18226 ( .A(n9334), .Z(n184) );
  HS65_LS_IVX2 U18227 ( .A(n9340), .Z(n653) );
  HS65_LS_IVX2 U18228 ( .A(n9355), .Z(n429) );
  HS65_LS_IVX2 U18229 ( .A(n9313), .Z(n116) );
  HS65_LS_IVX2 U18230 ( .A(n9329), .Z(n603) );
  HS65_LS_IVX2 U18231 ( .A(n9366), .Z(n209) );
  HS65_LS_IVX2 U18232 ( .A(sa03[2]), .Z(n183) );
  HS65_LS_AO22X4 U18233 ( .A(key[22]), .B(n9856), .C(n1037), .D(n9864), .Z(
        w3[22]) );
  HS65_LSS_XOR2X3 U18234 ( .A(n892), .B(n1038), .Z(n1037) );
  HS65_LS_AO22X4 U18235 ( .A(key[5]), .B(n9857), .C(n1071), .D(n9865), .Z(
        w3[5]) );
  HS65_LSS_XOR2X3 U18236 ( .A(n809), .B(n1072), .Z(n1071) );
  HS65_LS_OAI22X1 U18237 ( .A(n5978), .B(n9145), .C(n9137), .D(n5979), .Z(
        sa01[0]) );
  HS65_LSS_XNOR2X3 U18238 ( .A(n9234), .B(n9677), .Z(n5978) );
  HS65_LSS_XOR3X2 U18239 ( .A(n274), .B(n5980), .C(n5981), .Z(n5979) );
  HS65_LSS_XOR2X3 U18240 ( .A(n9234), .B(n2769), .Z(n5981) );
  HS65_LS_OAI22X1 U18241 ( .A(n9477), .B(n9582), .C(n9586), .D(n9422), .Z(
        sa12[6]) );
  HS65_LSS_XNOR2X3 U18242 ( .A(n9250), .B(n9643), .Z(n7576) );
  HS65_LSS_XOR3X2 U18243 ( .A(n7550), .B(n7578), .C(n7579), .Z(n7577) );
  HS65_LSS_XOR2X3 U18244 ( .A(n9250), .B(n2791), .Z(n7579) );
  HS65_LS_OAI22X1 U18245 ( .A(n2631), .B(n9145), .C(n9138), .D(n2632), .Z(
        sa32[0]) );
  HS65_LSS_XNOR2X3 U18246 ( .A(n9282), .B(n9621), .Z(n2631) );
  HS65_LSS_XOR3X2 U18247 ( .A(n2626), .B(n2633), .C(n2634), .Z(n2632) );
  HS65_LSS_XOR2X3 U18248 ( .A(n9282), .B(n316), .Z(n2634) );
  HS65_LS_OAI22X1 U18249 ( .A(n7573), .B(n9142), .C(n9139), .D(n7574), .Z(
        sa12[7]) );
  HS65_LSS_XNOR2X3 U18250 ( .A(n9280), .B(n9644), .Z(n7573) );
  HS65_LSS_XOR3X2 U18251 ( .A(n7542), .B(n7545), .C(n7575), .Z(n7574) );
  HS65_LSS_XOR2X3 U18252 ( .A(n9280), .B(n317), .Z(n7575) );
  HS65_LS_OAI22X1 U18253 ( .A(n5985), .B(n9142), .C(n9137), .D(n5986), .Z(
        sa11[6]) );
  HS65_LSS_XNOR2X3 U18254 ( .A(n9233), .B(n9675), .Z(n5985) );
  HS65_LSS_XOR3X2 U18255 ( .A(n5958), .B(n5987), .C(n5988), .Z(n5986) );
  HS65_LSS_XOR2X3 U18256 ( .A(n9233), .B(n52), .Z(n5988) );
  HS65_LS_OAI22X1 U18257 ( .A(n4392), .B(n9147), .C(n9140), .D(n4393), .Z(
        sa10[6]) );
  HS65_LSS_XNOR2X3 U18258 ( .A(n9271), .B(n9707), .Z(n4392) );
  HS65_LSS_XOR3X2 U18259 ( .A(n4365), .B(n4394), .C(n4395), .Z(n4393) );
  HS65_LSS_XOR2X3 U18260 ( .A(n9271), .B(n232), .Z(n4395) );
  HS65_LS_OAI22X1 U18261 ( .A(n8032), .B(n9147), .C(n9137), .D(n8033), .Z(
        sa32[5]) );
  HS65_LSS_XNOR2X3 U18262 ( .A(n9287), .B(n9626), .Z(n8032) );
  HS65_LSS_XOR3X2 U18263 ( .A(n7550), .B(n7588), .C(n8034), .Z(n8033) );
  HS65_LSS_XOR2X3 U18264 ( .A(n9287), .B(n3013), .Z(n8034) );
  HS65_LS_AO22X4 U18265 ( .A(key[23]), .B(n9856), .C(n1035), .D(n9864), .Z(
        w3[23]) );
  HS65_LSS_XOR2X3 U18266 ( .A(n893), .B(n1036), .Z(n1035) );
  HS65_LS_IVX2 U18267 ( .A(n9399), .Z(n604) );
  HS65_LS_IVX2 U18268 ( .A(n9309), .Z(n117) );
  HS65_LS_IVX2 U18269 ( .A(n9403), .Z(n333) );
  HS65_LS_IVX2 U18270 ( .A(n9357), .Z(n339) );
  HS65_LS_IVX2 U18271 ( .A(n9382), .Z(n382) );
  HS65_LS_IVX2 U18272 ( .A(n9375), .Z(n384) );
  HS65_LS_IVX2 U18273 ( .A(n9342), .Z(n621) );
  HS65_LS_IVX2 U18274 ( .A(n9344), .Z(n360) );
  HS65_LS_IVX2 U18275 ( .A(n9354), .Z(n490) );
  HS65_LS_IVX2 U18276 ( .A(n9352), .Z(n271) );
  HS65_LS_IVX2 U18277 ( .A(n9321), .Z(n708) );
  HS65_LS_IVX2 U18278 ( .A(sa33[3]), .Z(n44) );
  HS65_LS_IVX2 U18279 ( .A(n9343), .Z(n418) );
  HS65_LS_IVX2 U18280 ( .A(n9350), .Z(n449) );
  HS65_LS_IVX2 U18281 ( .A(n9327), .Z(n672) );
  HS65_LS_IVX2 U18282 ( .A(n9383), .Z(n642) );
  HS65_LS_IVX2 U18283 ( .A(sa32[7]), .Z(n206) );
  HS65_LS_IVX2 U18284 ( .A(n9315), .Z(n163) );
  HS65_LS_IVX2 U18285 ( .A(n9299), .Z(n161) );
  HS65_LS_IVX2 U18286 ( .A(n9247), .Z(n134) );
  HS65_LS_IVX2 U18287 ( .A(n9240), .Z(n313) );
  HS65_LS_IVX2 U18288 ( .A(sa23[3]), .Z(n92) );
  HS65_LS_IVX2 U18289 ( .A(n9237), .Z(n570) );
  HS65_LS_IVX2 U18290 ( .A(n9353), .Z(n526) );
  HS65_LS_IVX2 U18291 ( .A(n9360), .Z(n405) );
  HS65_LS_IVX2 U18292 ( .A(sa32[1]), .Z(n229) );
  HS65_LS_OAI22X1 U18293 ( .A(n5982), .B(n9146), .C(n9137), .D(n5983), .Z(
        sa11[7]) );
  HS65_LSS_XNOR2X3 U18294 ( .A(n9231), .B(n9676), .Z(n5982) );
  HS65_LSS_XOR3X2 U18295 ( .A(n5950), .B(n5954), .C(n5984), .Z(n5983) );
  HS65_LSS_XNOR2X3 U18296 ( .A(n9231), .B(n3219), .Z(n5984) );
  HS65_LS_OAI22X1 U18297 ( .A(n4446), .B(n9147), .C(n9138), .D(n4447), .Z(
        sa20[0]) );
  HS65_LSS_XNOR2X3 U18298 ( .A(n9258), .B(n9693), .Z(n4446) );
  HS65_LSS_XOR3X2 U18299 ( .A(n4357), .B(n4419), .C(n4448), .Z(n4447) );
  HS65_LSS_XNOR2X3 U18300 ( .A(n9258), .B(n2825), .Z(n4448) );
  HS65_LS_OAI22X1 U18301 ( .A(n4389), .B(n9147), .C(n9141), .D(n4390), .Z(
        sa10[7]) );
  HS65_LSS_XNOR2X3 U18302 ( .A(n9261), .B(n9708), .Z(n4389) );
  HS65_LSS_XOR3X2 U18303 ( .A(n4357), .B(n4361), .C(n4391), .Z(n4390) );
  HS65_LSS_XNOR2X3 U18304 ( .A(n9261), .B(n3544), .Z(n4391) );
  HS65_LS_OAI22X1 U18305 ( .A(n6042), .B(n9147), .C(n9136), .D(n6043), .Z(
        sa31[7]) );
  HS65_LSS_XNOR2X3 U18306 ( .A(n9229), .B(n9660), .Z(n6042) );
  HS65_LSS_XOR3X2 U18307 ( .A(n274), .B(n5987), .C(n6044), .Z(n6043) );
  HS65_LSS_XNOR2X3 U18308 ( .A(n9229), .B(n2800), .Z(n6044) );
  HS65_LS_OAI22X1 U18309 ( .A(n4449), .B(n9146), .C(n9138), .D(n4450), .Z(
        sa30[7]) );
  HS65_LSS_XNOR2X3 U18310 ( .A(n9263), .B(n9692), .Z(n4449) );
  HS65_LSS_XOR3X2 U18311 ( .A(n451), .B(n4394), .C(n4451), .Z(n4450) );
  HS65_LSS_XNOR2X3 U18312 ( .A(n9263), .B(n2808), .Z(n4451) );
  HS65_LS_OAI22X1 U18313 ( .A(n6010), .B(n9147), .C(n9136), .D(n6011), .Z(
        sa11[0]) );
  HS65_LSS_XNOR2X3 U18314 ( .A(n9230), .B(n9669), .Z(n6010) );
  HS65_LSS_XOR3X2 U18315 ( .A(n5995), .B(n6012), .C(n6013), .Z(n6011) );
  HS65_LSS_XNOR2X3 U18316 ( .A(n9230), .B(n2793), .Z(n6013) );
  HS65_LS_OAI22X1 U18317 ( .A(n7711), .B(n9145), .C(n9137), .D(n7712), .Z(
        sa22[0]) );
  HS65_LSS_XNOR2X3 U18318 ( .A(n9297), .B(n9629), .Z(n7711) );
  HS65_LSS_XOR3X2 U18319 ( .A(n2629), .B(n7542), .C(n7713), .Z(n7712) );
  HS65_LSS_XNOR2X3 U18320 ( .A(n9297), .B(n2809), .Z(n7713) );
  HS65_LS_OAI22X1 U18321 ( .A(n6039), .B(n9147), .C(n9136), .D(n6040), .Z(
        sa21[0]) );
  HS65_LSS_XNOR2X3 U18322 ( .A(n9232), .B(n9661), .Z(n6039) );
  HS65_LSS_XOR3X2 U18323 ( .A(n5950), .B(n6012), .C(n6041), .Z(n6040) );
  HS65_LSS_XNOR2X3 U18324 ( .A(n9232), .B(n2817), .Z(n6041) );
  HS65_LS_OAI22X1 U18325 ( .A(n8852), .B(n9146), .C(n9136), .D(n8853), .Z(
        sa32[2]) );
  HS65_LSS_XNOR2X3 U18326 ( .A(n9292), .B(n9623), .Z(n8852) );
  HS65_LSS_XOR3X2 U18327 ( .A(n7565), .B(n7600), .C(n8854), .Z(n8853) );
  HS65_LSS_XNOR2X3 U18328 ( .A(n9292), .B(n3010), .Z(n8854) );
  HS65_LS_OAI22X1 U18329 ( .A(n7085), .B(n9148), .C(n9138), .D(n7086), .Z(
        sa31[2]) );
  HS65_LSS_XNOR2X3 U18330 ( .A(n9213), .B(n9655), .Z(n7085) );
  HS65_LSS_XOR3X2 U18331 ( .A(n5972), .B(n6009), .C(n7087), .Z(n7086) );
  HS65_LSS_XNOR2X3 U18332 ( .A(n9213), .B(n3018), .Z(n7087) );
  HS65_LS_OAI22X1 U18333 ( .A(n6214), .B(n9148), .C(n9141), .D(n6215), .Z(
        sa31[5]) );
  HS65_LSS_XNOR2X3 U18334 ( .A(n9212), .B(n9658), .Z(n6214) );
  HS65_LSS_XOR3X2 U18335 ( .A(n5958), .B(n5997), .C(n6216), .Z(n6215) );
  HS65_LSS_XNOR2X3 U18336 ( .A(n9212), .B(n3217), .Z(n6216) );
  HS65_LS_OAI22X1 U18337 ( .A(n4524), .B(n9147), .C(n9138), .D(n4525), .Z(
        sa30[6]) );
  HS65_LSS_XNOR2X3 U18338 ( .A(n9268), .B(n9691), .Z(n4524) );
  HS65_LSS_XOR3X2 U18339 ( .A(n4361), .B(n4398), .C(n4526), .Z(n4525) );
  HS65_LSS_XNOR2X3 U18340 ( .A(n9268), .B(n3543), .Z(n4526) );
  HS65_LS_OAI22X1 U18341 ( .A(n6117), .B(n9147), .C(n9136), .D(n6118), .Z(
        sa31[6]) );
  HS65_LSS_XNOR2X3 U18342 ( .A(n9227), .B(n9659), .Z(n6117) );
  HS65_LSS_XOR3X2 U18343 ( .A(n5954), .B(n5991), .C(n6119), .Z(n6118) );
  HS65_LSS_XNOR2X3 U18344 ( .A(n9227), .B(n3218), .Z(n6119) );
  HS65_LS_OAI22X1 U18345 ( .A(n5675), .B(n9148), .C(n9138), .D(n5676), .Z(
        sa30[0]) );
  HS65_LSS_XNOR2X3 U18346 ( .A(n9257), .B(n9685), .Z(n5675) );
  HS65_LSS_XOR3X2 U18347 ( .A(n4387), .B(n4813), .C(n5677), .Z(n5676) );
  HS65_LSS_XNOR2X3 U18348 ( .A(n9257), .B(n3220), .Z(n5677) );
  HS65_LS_OAI22X1 U18349 ( .A(n7267), .B(n9148), .C(n9137), .D(n7268), .Z(
        sa31[0]) );
  HS65_LSS_XNOR2X3 U18350 ( .A(n9228), .B(n9653), .Z(n7267) );
  HS65_LSS_XOR3X2 U18351 ( .A(n5980), .B(n6406), .C(n7269), .Z(n7268) );
  HS65_LSS_XNOR2X3 U18352 ( .A(n9228), .B(n3016), .Z(n7269) );
  HS65_LS_OAI22X1 U18353 ( .A(n7570), .B(n9142), .C(n9138), .D(n7571), .Z(
        sa02[0]) );
  HS65_LSS_XNOR2X3 U18354 ( .A(n9281), .B(n9645), .Z(n7570) );
  HS65_LSS_XNOR3X2 U18355 ( .A(n7556), .B(n2633), .C(n7572), .Z(n7571) );
  HS65_LSS_XNOR2X3 U18356 ( .A(n2761), .B(n9281), .Z(n7572) );
  HS65_LS_OAI22X1 U18357 ( .A(n5493), .B(n9145), .C(n9138), .D(n5494), .Z(
        sa30[2]) );
  HS65_LSS_XNOR2X3 U18358 ( .A(n9225), .B(n9687), .Z(n5493) );
  HS65_LSS_XOR3X2 U18359 ( .A(n4379), .B(n4416), .C(n5495), .Z(n5494) );
  HS65_LSS_XNOR2X3 U18360 ( .A(n9225), .B(n3222), .Z(n5495) );
  HS65_LS_OAI22X1 U18361 ( .A(n7941), .B(n9145), .C(n9138), .D(n7942), .Z(
        sa32[6]) );
  HS65_LSS_XNOR2X3 U18362 ( .A(n9291), .B(n9627), .Z(n7941) );
  HS65_LSS_XOR3X2 U18363 ( .A(n7582), .B(n7545), .C(n7943), .Z(n7942) );
  HS65_LSS_XOR2X3 U18364 ( .A(n3014), .B(n9291), .Z(n7943) );
  HS65_LS_OAI22X1 U18365 ( .A(n4621), .B(n9148), .C(n9138), .D(n4622), .Z(
        sa30[5]) );
  HS65_LSS_XNOR2X3 U18366 ( .A(n9226), .B(n9690), .Z(n4621) );
  HS65_LSS_XOR3X2 U18367 ( .A(n4365), .B(n4404), .C(n4623), .Z(n4622) );
  HS65_LSS_XNOR2X3 U18368 ( .A(n9226), .B(n3225), .Z(n4623) );
  HS65_LS_OAI22X1 U18369 ( .A(n8201), .B(n9145), .C(n9136), .D(n8202), .Z(
        sa32[4]) );
  HS65_LSS_XNOR2X3 U18370 ( .A(n9289), .B(n9625), .Z(n8201) );
  HS65_LSS_XOR3X2 U18371 ( .A(n7554), .B(n8203), .C(n7592), .Z(n8202) );
  HS65_LSS_XOR3X2 U18372 ( .A(n9289), .B(n2626), .C(n3012), .Z(n8203) );
  HS65_LS_OAI22X1 U18373 ( .A(n6018), .B(n9147), .C(n9136), .D(n6019), .Z(
        sa21[6]) );
  HS65_LSS_XNOR2X3 U18374 ( .A(n9224), .B(n9667), .Z(n6018) );
  HS65_LSS_XOR3X2 U18375 ( .A(n2823), .B(n5987), .C(n6020), .Z(n6019) );
  HS65_LSS_XOR3X2 U18376 ( .A(n2774), .B(n9224), .C(n2798), .Z(n6020) );
  HS65_LS_OAI22X1 U18377 ( .A(n7610), .B(n9142), .C(n9138), .D(n7611), .Z(
        sa22[5]) );
  HS65_LSS_XNOR2X3 U18378 ( .A(n9286), .B(n9634), .Z(n7610) );
  HS65_LSS_XOR3X2 U18379 ( .A(n2814), .B(n7612), .C(n7582), .Z(n7611) );
  HS65_LSS_XOR3X2 U18380 ( .A(n2765), .B(n9286), .C(n2789), .Z(n7612) );
  HS65_LS_OAI22X1 U18381 ( .A(n7621), .B(n9147), .C(n9140), .D(n7622), .Z(
        sa22[2]) );
  HS65_LSS_XNOR2X3 U18382 ( .A(n9295), .B(n9631), .Z(n7621) );
  HS65_LSS_XOR3X2 U18383 ( .A(n2811), .B(n7623), .C(n7595), .Z(n7622) );
  HS65_LSS_XOR3X2 U18384 ( .A(n2786), .B(n9295), .C(n2762), .Z(n7623) );
  HS65_LS_OAI22X1 U18385 ( .A(n7613), .B(n9142), .C(n9141), .D(n7614), .Z(
        sa22[4]) );
  HS65_LSS_XNOR2X3 U18386 ( .A(n9288), .B(n9633), .Z(n7613) );
  HS65_LSS_XOR3X2 U18387 ( .A(n7588), .B(n7615), .C(n7616), .Z(n7614) );
  HS65_LSS_XOR3X2 U18388 ( .A(n2764), .B(n9288), .C(n2788), .Z(n7616) );
  HS65_LS_OAI22X1 U18389 ( .A(n8490), .B(n9145), .C(n9137), .D(n8491), .Z(
        sa32[3]) );
  HS65_LSS_XNOR2X3 U18390 ( .A(n9296), .B(n9624), .Z(n8490) );
  HS65_LSS_XOR3X2 U18391 ( .A(n7560), .B(n8492), .C(n7595), .Z(n8491) );
  HS65_LSS_XNOR3X2 U18392 ( .A(n9296), .B(n2626), .C(n3011), .Z(n8492) );
  HS65_LS_OAI22X1 U18393 ( .A(n7163), .B(n9145), .C(n9137), .D(n7164), .Z(
        sa31[1]) );
  HS65_LSS_XNOR2X3 U18394 ( .A(n9223), .B(n9654), .Z(n7163) );
  HS65_LSS_XOR3X2 U18395 ( .A(n6012), .B(n7165), .C(n6406), .Z(n7164) );
  HS65_LSS_XNOR3X2 U18396 ( .A(n9223), .B(n5975), .C(n3017), .Z(n7165) );
  HS65_LS_OAI22X1 U18397 ( .A(n6021), .B(n9146), .C(n9136), .D(n6022), .Z(
        sa21[5]) );
  HS65_LSS_XNOR2X3 U18398 ( .A(n9209), .B(n9666), .Z(n6021) );
  HS65_LSS_XNOR3X2 U18399 ( .A(n2822), .B(n6023), .C(n5991), .Z(n6022) );
  HS65_LSS_XOR3X2 U18400 ( .A(n2773), .B(n9209), .C(n2797), .Z(n6023) );
  HS65_LS_OAI22X1 U18401 ( .A(n6032), .B(n9148), .C(n9136), .D(n6033), .Z(
        sa21[2]) );
  HS65_LSS_XNOR2X3 U18402 ( .A(n9210), .B(n9663), .Z(n6032) );
  HS65_LSS_XOR3X2 U18403 ( .A(n2819), .B(n6034), .C(n6004), .Z(n6033) );
  HS65_LSS_XOR3X2 U18404 ( .A(n2770), .B(n9210), .C(n2794), .Z(n6034) );
  HS65_LS_OAI22X1 U18405 ( .A(n7547), .B(n9142), .C(n9136), .D(n7548), .Z(
        sa02[5]) );
  HS65_LSS_XNOR2X3 U18406 ( .A(n9275), .B(n9650), .Z(n7547) );
  HS65_LSS_XOR3X2 U18407 ( .A(n3012), .B(n7549), .C(n7550), .Z(n7548) );
  HS65_LSS_XOR3X2 U18408 ( .A(n2766), .B(n9275), .C(n2813), .Z(n7549) );
  HS65_LS_OAI22X1 U18409 ( .A(n7551), .B(n9142), .C(n9136), .D(n7552), .Z(
        sa02[4]) );
  HS65_LSS_XNOR2X3 U18410 ( .A(n9276), .B(n9649), .Z(n7551) );
  HS65_LSS_XOR3X2 U18411 ( .A(n7553), .B(n7554), .C(n7555), .Z(n7552) );
  HS65_LSS_XOR3X2 U18412 ( .A(n9276), .B(n364), .C(n2812), .Z(n7555) );
  HS65_LS_OAI22X1 U18413 ( .A(n6024), .B(n9145), .C(n9136), .D(n6025), .Z(
        sa21[4]) );
  HS65_LSS_XNOR2X3 U18414 ( .A(n9208), .B(n9665), .Z(n6024) );
  HS65_LSS_XOR3X2 U18415 ( .A(n5997), .B(n6026), .C(n6027), .Z(n6025) );
  HS65_LSS_XOR3X2 U18416 ( .A(n2772), .B(n9208), .C(n2796), .Z(n6027) );
  HS65_LS_OAI22X1 U18417 ( .A(n9476), .B(n9576), .C(n9586), .D(n9421), .Z(
        sa32[1]) );
  HS65_LSS_XNOR2X3 U18418 ( .A(n9285), .B(n9622), .Z(n2624) );
  HS65_LSS_XOR3X2 U18419 ( .A(n2626), .B(n2627), .C(n2628), .Z(n2625) );
  HS65_LSS_XOR3X2 U18420 ( .A(n9285), .B(n2629), .C(n2630), .Z(n2627) );
  HS65_LS_OAI22X1 U18421 ( .A(n5998), .B(n9145), .C(n9137), .D(n5999), .Z(
        sa11[3]) );
  HS65_LSS_XNOR2X3 U18422 ( .A(n9218), .B(n9672), .Z(n5998) );
  HS65_LSS_XOR3X2 U18423 ( .A(n5995), .B(n6000), .C(n6001), .Z(n5999) );
  HS65_LSS_XOR3X2 U18424 ( .A(n9218), .B(n5972), .C(n2796), .Z(n6000) );
  HS65_LS_OAI22X1 U18425 ( .A(n5964), .B(n9146), .C(n9137), .D(n5965), .Z(
        sa01[3]) );
  HS65_LSS_XNOR2X3 U18426 ( .A(n9220), .B(n9680), .Z(n5964) );
  HS65_LSS_XOR3X2 U18427 ( .A(n5966), .B(n5967), .C(n5968), .Z(n5965) );
  HS65_LSS_XOR3X2 U18428 ( .A(n9220), .B(n2772), .C(n2819), .Z(n5968) );
  HS65_LS_OAI22X1 U18429 ( .A(n7617), .B(n9147), .C(n9136), .D(n7618), .Z(
        sa22[3]) );
  HS65_LSS_XNOR2X3 U18430 ( .A(n9290), .B(n9632), .Z(n7617) );
  HS65_LSS_XOR3X2 U18431 ( .A(n7619), .B(n7592), .C(n7620), .Z(n7618) );
  HS65_LSS_XOR3X2 U18432 ( .A(n9290), .B(n2763), .C(n577), .Z(n7620) );
  HS65_LS_OAI22X1 U18433 ( .A(n7648), .B(n9147), .C(n9140), .D(n7649), .Z(
        sa22[1]) );
  HS65_LSS_XNOR2X3 U18434 ( .A(n9293), .B(n9630), .Z(n7648) );
  HS65_LSS_XOR3X2 U18435 ( .A(n7650), .B(n7600), .C(n7651), .Z(n7649) );
  HS65_LSS_XOR3X2 U18436 ( .A(n9293), .B(n2810), .C(n2761), .Z(n7651) );
  HS65_LS_OAI22X1 U18437 ( .A(n9475), .B(n9576), .C(n9584), .D(n9420), .Z(
        sa20[1]) );
  HS65_LSS_XNOR2X3 U18438 ( .A(n9264), .B(n9694), .Z(n4442) );
  HS65_LSS_XOR3X2 U18439 ( .A(n4444), .B(n4416), .C(n4445), .Z(n4443) );
  HS65_LSS_XOR2X3 U18440 ( .A(n2826), .B(n4357), .Z(n4444) );
  HS65_LS_OAI22X1 U18441 ( .A(n6035), .B(n9147), .C(n9136), .D(n6036), .Z(
        sa21[1]) );
  HS65_LSS_XNOR2X3 U18442 ( .A(n9221), .B(n9662), .Z(n6035) );
  HS65_LSS_XOR3X2 U18443 ( .A(n6037), .B(n6009), .C(n6038), .Z(n6036) );
  HS65_LSS_XOR2X3 U18444 ( .A(n2818), .B(n5950), .Z(n6037) );
  HS65_LS_OAI22X1 U18445 ( .A(n6006), .B(n9145), .C(n9136), .D(n6007), .Z(
        sa11[1]) );
  HS65_LSS_XNOR2X3 U18446 ( .A(n9219), .B(n9670), .Z(n6006) );
  HS65_LSS_XOR3X2 U18447 ( .A(n5995), .B(n6008), .C(n6009), .Z(n6007) );
  HS65_LSS_XOR3X2 U18448 ( .A(n9219), .B(n5980), .C(n51), .Z(n6008) );
  HS65_LS_OAI22X1 U18449 ( .A(n6403), .B(n9146), .C(n9137), .D(n6404), .Z(
        sa31[4]) );
  HS65_LSS_XNOR2X3 U18450 ( .A(n9207), .B(n9657), .Z(n6403) );
  HS65_LSS_XOR3X2 U18451 ( .A(n6001), .B(n6405), .C(n6406), .Z(n6404) );
  HS65_LSS_XNOR3X2 U18452 ( .A(n9207), .B(n5962), .C(n3216), .Z(n6405) );
  HS65_LS_OAI22X1 U18453 ( .A(n4431), .B(n9145), .C(n9139), .D(n4432), .Z(
        sa20[4]) );
  HS65_LSS_XNOR2X3 U18454 ( .A(n9214), .B(n9697), .Z(n4431) );
  HS65_LSS_XOR3X2 U18455 ( .A(n4404), .B(n4433), .C(n4434), .Z(n4432) );
  HS65_LSS_XOR3X2 U18456 ( .A(n2780), .B(n9214), .C(n2804), .Z(n4434) );
  HS65_LS_OAI22X1 U18457 ( .A(n5993), .B(n9145), .C(n9137), .D(n5994), .Z(
        sa11[4]) );
  HS65_LSS_XNOR2X3 U18458 ( .A(n9206), .B(n9673), .Z(n5993) );
  HS65_LSS_XOR3X2 U18459 ( .A(n5995), .B(n5996), .C(n5997), .Z(n5994) );
  HS65_LSS_XOR3X2 U18460 ( .A(n9206), .B(n5967), .C(n2797), .Z(n5996) );
  HS65_LS_OAI22X1 U18461 ( .A(n7584), .B(n9142), .C(n9140), .D(n7585), .Z(
        sa12[4]) );
  HS65_LSS_XNOR2X3 U18462 ( .A(n9251), .B(n9641), .Z(n7584) );
  HS65_LSS_XOR3X2 U18463 ( .A(n7586), .B(n7587), .C(n7588), .Z(n7585) );
  HS65_LSS_XOR3X2 U18464 ( .A(n9251), .B(n7560), .C(n2789), .Z(n7587) );
  HS65_LS_OAI22X1 U18465 ( .A(n9474), .B(n9582), .C(n9584), .D(n9419), .Z(
        sa22[7]) );
  HS65_LSS_XNOR2X3 U18466 ( .A(n9254), .B(n9636), .Z(n7604) );
  HS65_LSS_XOR3X2 U18467 ( .A(n2791), .B(n7606), .C(n7556), .Z(n7605) );
  HS65_LSS_XNOR3X2 U18468 ( .A(n2768), .B(n9254), .C(n2767), .Z(n7606) );
  HS65_LS_OAI22X1 U18469 ( .A(n7566), .B(n9142), .C(n9140), .D(n7567), .Z(
        sa02[1]) );
  HS65_LSS_XNOR2X3 U18470 ( .A(n9279), .B(n9646), .Z(n7566) );
  HS65_LSS_XOR2X3 U18471 ( .A(n7568), .B(n7569), .Z(n7567) );
  HS65_LSS_XOR3X2 U18472 ( .A(n9279), .B(n316), .C(n2809), .Z(n7568) );
  HS65_LS_OAI22X1 U18473 ( .A(n6014), .B(n9146), .C(n9136), .D(n6015), .Z(
        sa21[7]) );
  HS65_LSS_XNOR2X3 U18474 ( .A(n9217), .B(n9668), .Z(n6014) );
  HS65_LSS_XOR3X2 U18475 ( .A(n2799), .B(n6016), .C(n6017), .Z(n6015) );
  HS65_LSS_XNOR3X2 U18476 ( .A(n2775), .B(n9217), .C(n2776), .Z(n6016) );
  HS65_LS_OAI22X1 U18477 ( .A(n4435), .B(n9148), .C(n9139), .D(n4436), .Z(
        sa20[3]) );
  HS65_LSS_XNOR2X3 U18478 ( .A(n9269), .B(n9696), .Z(n4435) );
  HS65_LSS_XOR3X2 U18479 ( .A(n4437), .B(n4408), .C(n4438), .Z(n4436) );
  HS65_LSS_XOR3X2 U18480 ( .A(n9269), .B(n2779), .C(n233), .Z(n4438) );
  HS65_LS_OAI22X1 U18481 ( .A(n6028), .B(n9148), .C(n9136), .D(n6029), .Z(
        sa21[3]) );
  HS65_LSS_XNOR2X3 U18482 ( .A(n9216), .B(n9664), .Z(n6028) );
  HS65_LSS_XOR3X2 U18483 ( .A(n6030), .B(n6001), .C(n6031), .Z(n6029) );
  HS65_LSS_XOR3X2 U18484 ( .A(n9216), .B(n2771), .C(n53), .Z(n6031) );
  HS65_LS_OAI22X1 U18485 ( .A(n4400), .B(n9147), .C(n9139), .D(n4401), .Z(
        sa10[4]) );
  HS65_LSS_XNOR2X3 U18486 ( .A(n9211), .B(n9705), .Z(n4400) );
  HS65_LSS_XOR3X2 U18487 ( .A(n4402), .B(n4403), .C(n4404), .Z(n4401) );
  HS65_LSS_XOR3X2 U18488 ( .A(n9211), .B(n4374), .C(n2805), .Z(n4403) );
  HS65_LSS_XOR2X3 U18489 ( .A(n2807), .B(n9273), .Z(n9735) );
  HS65_LSS_XOR2X3 U18490 ( .A(n3221), .B(n9262), .Z(n9724) );
  HS65_LSS_XOR2X3 U18491 ( .A(n3225), .B(n9194), .Z(n9720) );
  HS65_LSS_XOR2X3 U18492 ( .A(n3222), .B(n9192), .Z(n9723) );
  HS65_LSS_XOR2X3 U18493 ( .A(n3217), .B(n9200), .Z(n9752) );
  HS65_LSS_XOR2X3 U18494 ( .A(n3544), .B(n9248), .Z(n9718) );
  HS65_LSS_XOR2X3 U18495 ( .A(n3018), .B(n9198), .Z(n9755) );
  HS65_LSS_XOR2X3 U18496 ( .A(n2803), .B(n9196), .Z(n9739) );
  HS65_LSS_XOR2X3 U18497 ( .A(n3224), .B(n9193), .Z(n9721) );
  HS65_LSS_XOR2X3 U18498 ( .A(n3223), .B(n9265), .Z(n9722) );
  HS65_LSS_XOR2X3 U18499 ( .A(n3216), .B(n9197), .Z(n9753) );
  HS65_LSS_XOR2X3 U18500 ( .A(n2828), .B(n9270), .Z(n9730) );
  HS65_LS_AO22X4 U18501 ( .A(key[13]), .B(n9857), .C(n1055), .D(n9865), .Z(
        w3[13]) );
  HS65_LSS_XOR2X3 U18502 ( .A(n850), .B(n1056), .Z(n1055) );
  HS65_LS_AO22X4 U18503 ( .A(key[15]), .B(n9857), .C(n1051), .D(n9859), .Z(
        w3[15]) );
  HS65_LSS_XOR2X3 U18504 ( .A(n852), .B(n1052), .Z(n1051) );
  HS65_LS_AO22X4 U18505 ( .A(key[25]), .B(n9856), .C(n1031), .D(n9864), .Z(
        w3[25]) );
  HS65_LSS_XOR2X3 U18506 ( .A(n912), .B(n1032), .Z(n1031) );
  HS65_LS_OAI22X1 U18507 ( .A(n7557), .B(n9142), .C(n9136), .D(n7558), .Z(
        sa02[3]) );
  HS65_LSS_XOR2X3 U18508 ( .A(n942), .B(n9648), .Z(n7557) );
  HS65_LSS_XNOR3X2 U18509 ( .A(n7559), .B(n7560), .C(n7561), .Z(n7558) );
  HS65_LSS_XOR3X2 U18510 ( .A(n942), .B(n2764), .C(n2811), .Z(n7561) );
  HS65_LS_OAI22X1 U18511 ( .A(n7580), .B(n9142), .C(n9141), .D(n7581), .Z(
        sa12[5]) );
  HS65_LSS_XOR2X3 U18512 ( .A(n940), .B(n9642), .Z(n7580) );
  HS65_LSS_XNOR3X2 U18513 ( .A(n7554), .B(n7582), .C(n7583), .Z(n7581) );
  HS65_LSS_XOR2X3 U18514 ( .A(n940), .B(n2790), .Z(n7583) );
  HS65_LS_OAI22X1 U18515 ( .A(n2675), .B(n9144), .C(n9141), .D(n2676), .Z(
        sa03[1]) );
  HS65_LSS_XOR2X3 U18516 ( .A(n912), .B(n9614), .Z(n2675) );
  HS65_LSS_XNOR3X2 U18517 ( .A(n2677), .B(n2678), .C(n2679), .Z(n2676) );
  HS65_LSS_XOR3X2 U18518 ( .A(n2681), .B(n9337), .C(n2682), .Z(n2678) );
  HS65_LS_OAI22X1 U18519 ( .A(n9461), .B(n9580), .C(n9587), .D(n9418), .Z(
        sa23[1]) );
  HS65_LSS_XOR2X3 U18520 ( .A(n830), .B(n9598), .Z(n2753) );
  HS65_LSS_XNOR3X2 U18521 ( .A(n2721), .B(n2755), .C(n2756), .Z(n2754) );
  HS65_LSS_XOR3X2 U18522 ( .A(n2757), .B(n9176), .C(n2687), .Z(n2755) );
  HS65_LS_OAI22X1 U18523 ( .A(n4380), .B(n9143), .C(n9588), .D(n4381), .Z(
        sa00[1]) );
  HS65_LSS_XOR2X3 U18524 ( .A(n964), .B(n9710), .Z(n4380) );
  HS65_LSS_XNOR3X2 U18525 ( .A(n4382), .B(n4383), .C(n4384), .Z(n4381) );
  HS65_LSS_XOR3X2 U18526 ( .A(n2778), .B(n9262), .C(n2825), .Z(n4383) );
  HS65_LS_OAI22X1 U18527 ( .A(n5973), .B(n9145), .C(n9137), .D(n5974), .Z(
        sa01[1]) );
  HS65_LSS_XOR2X3 U18528 ( .A(n946), .B(n9678), .Z(n5973) );
  HS65_LSS_XNOR3X2 U18529 ( .A(n5975), .B(n5976), .C(n5977), .Z(n5974) );
  HS65_LS_IVX2 U18530 ( .A(n9204), .Z(n946) );
  HS65_LSS_XOR2X3 U18531 ( .A(n953), .B(n2393), .Z(n1015) );
  HS65_LS_NAND4ABX3 U18532 ( .A(n2394), .B(n2395), .C(n2396), .D(n2397), .Z(
        n2393) );
  HS65_LS_MX41X4 U18533 ( .D0(n897), .S0(n921), .D1(n925), .S1(n909), .D2(n895), .S2(n916), .D3(n927), .S3(n2306), .Z(n2395) );
  HS65_LS_AOI212X2 U18534 ( .A(n910), .B(n2398), .C(n926), .D(n2375), .E(n2399), .Z(n2397) );
  HS65_LSS_XNOR2X3 U18535 ( .A(n9261), .B(n1491), .Z(n995) );
  HS65_LS_NAND4ABX3 U18536 ( .A(n1492), .B(n1493), .C(n1494), .D(n1495), .Z(
        n1491) );
  HS65_LS_OAI212X3 U18537 ( .A(n1503), .B(n1504), .C(n1505), .D(n1506), .E(
        n1507), .Z(n1493) );
  HS65_LS_NAND4ABX3 U18538 ( .A(n1513), .B(n1514), .C(n1515), .D(n1516), .Z(
        n1492) );
  HS65_LS_OAI22X1 U18539 ( .A(n720), .B(n9866), .C(n988), .D(n9848), .Z(w0[30]) );
  HS65_LS_IVX2 U18540 ( .A(key[126]), .Z(n720) );
  HS65_LSS_XOR3X2 U18541 ( .A(n1382), .B(n9404), .C(n965), .Z(n992) );
  HS65_LS_NOR4ABX2 U18542 ( .A(n1383), .B(n1384), .C(n1385), .D(n1386), .Z(
        n1382) );
  HS65_LS_CBI4I1X3 U18543 ( .A(n1201), .B(n1129), .C(n1155), .D(n1334), .Z(
        n1386) );
  HS65_LS_CBI4I6X2 U18544 ( .A(n860), .B(n1356), .C(n881), .D(n1405), .Z(n1383) );
  HS65_LS_OAI22X1 U18545 ( .A(n4417), .B(n9147), .C(n9139), .D(n4418), .Z(
        sa10[0]) );
  HS65_LSS_XOR2X3 U18546 ( .A(n958), .B(n9701), .Z(n4417) );
  HS65_LSS_XOR3X2 U18547 ( .A(n4402), .B(n4419), .C(n4420), .Z(n4418) );
  HS65_LSS_XOR2X3 U18548 ( .A(n958), .B(n2801), .Z(n4420) );
  HS65_LS_OAI22X1 U18549 ( .A(n4425), .B(n9148), .C(n9139), .D(n4426), .Z(
        sa20[6]) );
  HS65_LSS_XOR2X3 U18550 ( .A(n956), .B(n9699), .Z(n4425) );
  HS65_LSS_XOR3X2 U18551 ( .A(n2831), .B(n4394), .C(n4427), .Z(n4426) );
  HS65_LSS_XOR3X2 U18552 ( .A(n2782), .B(n9273), .C(n2806), .Z(n4427) );
  HS65_LS_OAI22X1 U18553 ( .A(n5959), .B(n9146), .C(n9137), .D(n5960), .Z(
        sa01[4]) );
  HS65_LSS_XOR2X3 U18554 ( .A(n948), .B(n9681), .Z(n5959) );
  HS65_LSS_XOR3X2 U18555 ( .A(n5961), .B(n5962), .C(n5963), .Z(n5960) );
  HS65_LSS_XOR3X2 U18556 ( .A(n9197), .B(n2773), .C(n2820), .Z(n5963) );
  HS65_LS_OAI22X1 U18557 ( .A(n4405), .B(n9148), .C(n9139), .D(n4406), .Z(
        sa10[3]) );
  HS65_LSS_XOR2X3 U18558 ( .A(n961), .B(n9704), .Z(n4405) );
  HS65_LSS_XOR3X2 U18559 ( .A(n4402), .B(n4407), .C(n4408), .Z(n4406) );
  HS65_LSS_XOR3X2 U18560 ( .A(n9270), .B(n4379), .C(n2804), .Z(n4407) );
  HS65_LS_OAI22X1 U18561 ( .A(n5989), .B(n9148), .C(n9137), .D(n5990), .Z(
        sa11[5]) );
  HS65_LSS_XOR2X3 U18562 ( .A(n945), .B(n9674), .Z(n5989) );
  HS65_LSS_XOR3X2 U18563 ( .A(n5962), .B(n5991), .C(n5992), .Z(n5990) );
  HS65_LSS_XOR2X3 U18564 ( .A(n945), .B(n2798), .Z(n5992) );
  HS65_LS_OAI22X1 U18565 ( .A(n6002), .B(n9146), .C(n9137), .D(n6003), .Z(
        sa11[2]) );
  HS65_LSS_XOR2X3 U18566 ( .A(n944), .B(n9671), .Z(n6002) );
  HS65_LSS_XOR3X2 U18567 ( .A(n6004), .B(n5975), .C(n6005), .Z(n6003) );
  HS65_LSS_XOR2X3 U18568 ( .A(n2795), .B(n9201), .Z(n6005) );
  HS65_LS_OAI22X1 U18569 ( .A(n4409), .B(n9148), .C(n9139), .D(n4410), .Z(
        sa10[2]) );
  HS65_LSS_XOR2X3 U18570 ( .A(n960), .B(n9703), .Z(n4409) );
  HS65_LSS_XOR3X2 U18571 ( .A(n4411), .B(n4382), .C(n4412), .Z(n4410) );
  HS65_LSS_XOR2X3 U18572 ( .A(n2803), .B(n9195), .Z(n4412) );
  HS65_LS_OAI22X1 U18573 ( .A(n4396), .B(n9148), .C(n9139), .D(n4397), .Z(
        sa10[5]) );
  HS65_LSS_XOR2X3 U18574 ( .A(n962), .B(n9706), .Z(n4396) );
  HS65_LSS_XOR3X2 U18575 ( .A(n4369), .B(n4398), .C(n4399), .Z(n4397) );
  HS65_LSS_XOR2X3 U18576 ( .A(n962), .B(n2806), .Z(n4399) );
  HS65_LS_OAI22X1 U18577 ( .A(n4439), .B(n9148), .C(n9139), .D(n4440), .Z(
        sa20[2]) );
  HS65_LSS_XOR2X3 U18578 ( .A(n955), .B(n9695), .Z(n4439) );
  HS65_LSS_XOR3X2 U18579 ( .A(n2827), .B(n4441), .C(n4411), .Z(n4440) );
  HS65_LSS_XOR3X2 U18580 ( .A(n2778), .B(n9196), .C(n2802), .Z(n4441) );
  HS65_LS_OAI22X1 U18581 ( .A(n4371), .B(n9143), .C(n9137), .D(n4372), .Z(
        sa00[3]) );
  HS65_LSS_XOR2X3 U18582 ( .A(n966), .B(n9712), .Z(n4371) );
  HS65_LSS_XOR3X2 U18583 ( .A(n4373), .B(n4374), .C(n4375), .Z(n4372) );
  HS65_LSS_XOR3X2 U18584 ( .A(n9265), .B(n2780), .C(n2827), .Z(n4375) );
  HS65_LS_OAI22X1 U18585 ( .A(n4366), .B(n9143), .C(n9136), .D(n4367), .Z(
        sa00[4]) );
  HS65_LSS_XOR2X3 U18586 ( .A(n967), .B(n9713), .Z(n4366) );
  HS65_LSS_XOR3X2 U18587 ( .A(n4368), .B(n4369), .C(n4370), .Z(n4367) );
  HS65_LSS_XOR3X2 U18588 ( .A(n9193), .B(n2781), .C(n2828), .Z(n4370) );
  HS65_LS_OAI22X1 U18589 ( .A(n2909), .B(n9143), .C(n9140), .D(n2910), .Z(
        sa33[6]) );
  HS65_LSS_XOR2X3 U18590 ( .A(n810), .B(n9595), .Z(n2909) );
  HS65_LSS_XOR3X2 U18591 ( .A(n2644), .B(n2699), .C(n2911), .Z(n2910) );
  HS65_LSS_XOR2X3 U18592 ( .A(n810), .B(n2640), .Z(n2911) );
  HS65_LS_OAI22X1 U18593 ( .A(n7601), .B(n9142), .C(n9141), .D(n7602), .Z(
        sa12[0]) );
  HS65_LSS_XOR2X3 U18594 ( .A(n936), .B(n9637), .Z(n7601) );
  HS65_LSS_XOR3X2 U18595 ( .A(n2629), .B(n7586), .C(n7603), .Z(n7602) );
  HS65_LSS_XOR2X3 U18596 ( .A(n936), .B(n2785), .Z(n7603) );
  HS65_LS_OAI22X1 U18597 ( .A(n2723), .B(n9144), .C(n9141), .D(n2724), .Z(
        sa13[0]) );
  HS65_LSS_XOR2X3 U18598 ( .A(n870), .B(n9605), .Z(n2723) );
  HS65_LSS_XOR3X2 U18599 ( .A(n2704), .B(n2725), .C(n2726), .Z(n2724) );
  HS65_LSS_XOR2X3 U18600 ( .A(n870), .B(n2727), .Z(n2726) );
  HS65_LS_OAI22X1 U18601 ( .A(n2683), .B(n9144), .C(n9141), .D(n2684), .Z(
        sa03[0]) );
  HS65_LSS_XOR2X3 U18602 ( .A(n911), .B(n9613), .Z(n2683) );
  HS65_LSS_XOR3X2 U18603 ( .A(n2661), .B(n2685), .C(n2686), .Z(n2684) );
  HS65_LSS_XOR2X3 U18604 ( .A(n911), .B(n2687), .Z(n2686) );
  HS65_LS_OAI22X1 U18605 ( .A(n2648), .B(n9144), .C(n9588), .D(n2649), .Z(
        sa03[5]) );
  HS65_LSS_XOR2X3 U18606 ( .A(n932), .B(n9618), .Z(n2648) );
  HS65_LSS_XOR3X2 U18607 ( .A(n630), .B(n2650), .C(n2651), .Z(n2649) );
  HS65_LSS_XOR3X2 U18608 ( .A(n2652), .B(n9181), .C(n2653), .Z(n2650) );
  HS65_LS_OAI22X1 U18609 ( .A(n2688), .B(n9144), .C(n9141), .D(n2689), .Z(
        sa13[7]) );
  HS65_LSS_XOR2X3 U18610 ( .A(n893), .B(n9612), .Z(n2688) );
  HS65_LSS_XOR3X2 U18611 ( .A(n2637), .B(n2644), .C(n2690), .Z(n2689) );
  HS65_LSS_XOR2X3 U18612 ( .A(n893), .B(n2691), .Z(n2690) );
  HS65_LS_OAI22X1 U18613 ( .A(n2692), .B(n9144), .C(n9141), .D(n2693), .Z(
        sa13[6]) );
  HS65_LSS_XOR2X3 U18614 ( .A(n892), .B(n9611), .Z(n2692) );
  HS65_LSS_XOR3X2 U18615 ( .A(n2651), .B(n2694), .C(n2695), .Z(n2693) );
  HS65_LSS_XOR2X3 U18616 ( .A(n892), .B(n2696), .Z(n2695) );
  HS65_LS_OAI22X1 U18617 ( .A(n9460), .B(n9581), .C(n9587), .D(n9417), .Z(
        sa23[4]) );
  HS65_LSS_XOR2X3 U18618 ( .A(n849), .B(n9601), .Z(n2741) );
  HS65_LSS_XOR3X2 U18619 ( .A(n2743), .B(n2706), .C(n2744), .Z(n2742) );
  HS65_LSS_XOR3X2 U18620 ( .A(n9185), .B(n630), .C(n2668), .Z(n2744) );
  HS65_LS_OAI22X1 U18621 ( .A(n4385), .B(n9143), .C(n9588), .D(n4386), .Z(
        sa00[0]) );
  HS65_LSS_XOR2X3 U18622 ( .A(n963), .B(n9709), .Z(n4385) );
  HS65_LSS_XOR3X2 U18623 ( .A(n451), .B(n4387), .C(n4388), .Z(n4386) );
  HS65_LSS_XOR2X3 U18624 ( .A(n9260), .B(n2777), .Z(n4388) );
  HS65_LS_OAI22X1 U18625 ( .A(n3020), .B(n9143), .C(n9140), .D(n3021), .Z(
        sa33[5]) );
  HS65_LSS_XOR2X3 U18626 ( .A(n809), .B(n9594), .Z(n3020) );
  HS65_LSS_XOR3X2 U18627 ( .A(n2651), .B(n2706), .C(n3022), .Z(n3021) );
  HS65_LSS_XOR2X3 U18628 ( .A(n809), .B(n2646), .Z(n3022) );
  HS65_LS_OAI22X1 U18629 ( .A(n2654), .B(n9144), .C(n9140), .D(n2655), .Z(
        sa03[4]) );
  HS65_LSS_XOR2X3 U18630 ( .A(n931), .B(n9617), .Z(n2654) );
  HS65_LSS_XOR3X2 U18631 ( .A(n2656), .B(n2657), .C(n2658), .Z(n2655) );
  HS65_LSS_XOR3X2 U18632 ( .A(n9179), .B(n187), .C(n2659), .Z(n2658) );
  HS65_LS_OAI22X1 U18633 ( .A(n2697), .B(n9144), .C(n9141), .D(n2698), .Z(
        sa13[5]) );
  HS65_LSS_XOR2X3 U18634 ( .A(n891), .B(n9610), .Z(n2697) );
  HS65_LSS_XOR3X2 U18635 ( .A(n2657), .B(n2699), .C(n2700), .Z(n2698) );
  HS65_LSS_XOR2X3 U18636 ( .A(n891), .B(n2701), .Z(n2700) );
  HS65_LS_OAI22X1 U18637 ( .A(n9459), .B(n9581), .C(n9585), .D(n9416), .Z(
        sa13[2]) );
  HS65_LSS_XOR2X3 U18638 ( .A(n872), .B(n9607), .Z(n2713) );
  HS65_LSS_XOR3X2 U18639 ( .A(n2677), .B(n2715), .C(n2716), .Z(n2714) );
  HS65_LSS_XOR2X3 U18640 ( .A(n872), .B(n2717), .Z(n2716) );
  HS65_LS_OAI22X1 U18641 ( .A(n2733), .B(n9144), .C(n9141), .D(n2734), .Z(
        sa23[6]) );
  HS65_LSS_XOR2X3 U18642 ( .A(n851), .B(n9603), .Z(n2733) );
  HS65_LSS_XOR3X2 U18643 ( .A(n186), .B(n2735), .C(n2694), .Z(n2734) );
  HS65_LSS_XOR3X2 U18644 ( .A(n851), .B(n409), .C(n2736), .Z(n2735) );
  HS65_LS_OAI22X1 U18645 ( .A(n3987), .B(n9143), .C(n9588), .D(n3988), .Z(
        sa33[1]) );
  HS65_LSS_XOR2X3 U18646 ( .A(n789), .B(n9590), .Z(n3987) );
  HS65_LSS_XOR3X2 U18647 ( .A(n2725), .B(n3989), .C(n3229), .Z(n3988) );
  HS65_LSS_XOR3X2 U18648 ( .A(n789), .B(n2677), .C(n2907), .Z(n3989) );
  HS65_LS_OAI22X1 U18649 ( .A(n9458), .B(n9581), .C(n9585), .D(n2671), .Z(
        sa03[2]) );
  HS65_LSS_XOR2X3 U18650 ( .A(n913), .B(n9615), .Z(n2670) );
  HS65_LSS_XOR3X2 U18651 ( .A(n9583), .B(n9415), .C(n9574), .Z(n2671) );
  HS65_LSS_XOR3X2 U18652 ( .A(n2674), .B(n9169), .C(n142), .Z(n2672) );
  HS65_LS_OAI22X1 U18653 ( .A(n3226), .B(n9143), .C(n9140), .D(n3227), .Z(
        sa33[4]) );
  HS65_LSS_XOR2X3 U18654 ( .A(n808), .B(n9593), .Z(n3226) );
  HS65_LSS_XOR3X2 U18655 ( .A(n2711), .B(n3228), .C(n3229), .Z(n3227) );
  HS65_LSS_XOR3X2 U18656 ( .A(n808), .B(n2657), .C(n2653), .Z(n3228) );
  HS65_LS_OAI22X1 U18657 ( .A(n2729), .B(n9144), .C(n9141), .D(n2730), .Z(
        sa23[7]) );
  HS65_LSS_XOR2X3 U18658 ( .A(n852), .B(n9604), .Z(n2729) );
  HS65_LSS_XOR3X2 U18659 ( .A(n188), .B(n2661), .C(n2731), .Z(n2730) );
  HS65_LSS_XOR3X2 U18660 ( .A(n2732), .B(n9338), .C(n2696), .Z(n2731) );
  HS65_LS_OAI22X1 U18661 ( .A(n9457), .B(n9581), .C(n9587), .D(n9456), .Z(
        sa03[3]) );
  HS65_LSS_XOR2X3 U18662 ( .A(n914), .B(n9616), .Z(n2662) );
  HS65_LSS_XOR2X3 U18663 ( .A(n2664), .B(n2665), .Z(n2663) );
  HS65_LSS_XOR3X2 U18664 ( .A(n914), .B(n141), .C(n2668), .Z(n2664) );
  HS65_LS_OAI22X1 U18665 ( .A(n9455), .B(n9581), .C(n9587), .D(n9454), .Z(
        sa23[3]) );
  HS65_LSS_XOR2X3 U18666 ( .A(n832), .B(n9600), .Z(n2746) );
  HS65_LSS_XOR2X3 U18667 ( .A(n2748), .B(n2749), .Z(n2747) );
  HS65_LSS_XOR3X2 U18668 ( .A(n832), .B(n408), .C(n2660), .Z(n2748) );
  HS65_LS_OAI22X1 U18669 ( .A(n3913), .B(n9143), .C(n9140), .D(n3914), .Z(
        sa33[2]) );
  HS65_LSS_XOR2X3 U18670 ( .A(n790), .B(n9591), .Z(n3913) );
  HS65_LSS_XOR3X2 U18671 ( .A(n2673), .B(n2721), .C(n3915), .Z(n3914) );
  HS65_LSS_XOR2X3 U18672 ( .A(n790), .B(n2669), .Z(n3915) );
  HS65_LS_OAI22X1 U18673 ( .A(n7593), .B(n9142), .C(n9139), .D(n7594), .Z(
        sa12[2]) );
  HS65_LSS_XOR2X3 U18674 ( .A(n938), .B(n9639), .Z(n7593) );
  HS65_LSS_XOR3X2 U18675 ( .A(n7595), .B(n2628), .C(n7596), .Z(n7594) );
  HS65_LSS_XOR2X3 U18676 ( .A(n2787), .B(n9255), .Z(n7596) );
  HS65_LS_OAI22X1 U18677 ( .A(n2833), .B(n9143), .C(n9140), .D(n2834), .Z(
        sa33[7]) );
  HS65_LSS_XOR2X3 U18678 ( .A(n811), .B(n9596), .Z(n2833) );
  HS65_LSS_XOR3X2 U18679 ( .A(n2661), .B(n2694), .C(n2835), .Z(n2834) );
  HS65_LSS_XOR2X3 U18680 ( .A(n811), .B(n2728), .Z(n2835) );
  HS65_LS_OAI22X1 U18681 ( .A(n2758), .B(n9143), .C(n9140), .D(n2759), .Z(
        sa23[0]) );
  HS65_LSS_XOR2X3 U18682 ( .A(n829), .B(n9597), .Z(n2758) );
  HS65_LSS_XOR3X2 U18683 ( .A(n2637), .B(n2725), .C(n2760), .Z(n2759) );
  HS65_LSS_XOR2X3 U18684 ( .A(n829), .B(n2680), .Z(n2760) );
  HS65_LS_OAI22X1 U18685 ( .A(n4081), .B(n9143), .C(n9588), .D(n4082), .Z(
        sa33[0]) );
  HS65_LSS_XOR2X3 U18686 ( .A(n788), .B(n9589), .Z(n4081) );
  HS65_LSS_XOR3X2 U18687 ( .A(n2685), .B(n3229), .C(n4083), .Z(n4082) );
  HS65_LSS_XOR2X3 U18688 ( .A(n788), .B(n2682), .Z(n4083) );
  HS65_LS_OAI22X1 U18689 ( .A(n2635), .B(n9145), .C(n9141), .D(n2636), .Z(
        sa03[7]) );
  HS65_LSS_XOR2X3 U18690 ( .A(n934), .B(n9620), .Z(n2635) );
  HS65_LSS_XOR3X2 U18691 ( .A(n631), .B(n2637), .C(n2638), .Z(n2636) );
  HS65_LSS_XOR3X2 U18692 ( .A(n2639), .B(n9183), .C(n2640), .Z(n2638) );
  HS65_LS_OAI22X1 U18693 ( .A(n2641), .B(n9145), .C(n9140), .D(n2642), .Z(
        sa03[6]) );
  HS65_LSS_XOR2X3 U18694 ( .A(n933), .B(n9619), .Z(n2641) );
  HS65_LSS_XOR3X2 U18695 ( .A(n632), .B(n2643), .C(n2644), .Z(n2642) );
  HS65_LS_IVX2 U18696 ( .A(n2647), .Z(n632) );
  HS65_LSS_XOR2X3 U18697 ( .A(n2781), .B(n954), .Z(n9745) );
  HS65_LS_OAI22X1 U18698 ( .A(n736), .B(n9861), .C(n1015), .D(n9854), .Z(
        \u0/N45 ) );
  HS65_LS_IVX2 U18699 ( .A(key[99]), .Z(n736) );
  HS65_LS_OAI22X1 U18700 ( .A(n762), .B(n9862), .C(n1066), .D(n9846), .Z(w2[8]) );
  HS65_LS_IVX2 U18701 ( .A(key[40]), .Z(n762) );
  HS65_LS_OAI22X1 U18702 ( .A(n767), .B(n9862), .C(n1076), .D(n9852), .Z(w2[3]) );
  HS65_LS_IVX2 U18703 ( .A(key[35]), .Z(n767) );
  HS65_LS_OAI22X1 U18704 ( .A(n760), .B(n9862), .C(n1062), .D(n9847), .Z(
        w2[10]) );
  HS65_LS_IVX2 U18705 ( .A(key[42]), .Z(n760) );
  HS65_LS_OAI22X1 U18706 ( .A(n763), .B(n9862), .C(n1068), .D(n9854), .Z(w2[7]) );
  HS65_LS_IVX2 U18707 ( .A(key[39]), .Z(n763) );
  HS65_LS_OAI22X1 U18708 ( .A(n761), .B(n9862), .C(n1064), .D(n9849), .Z(w2[9]) );
  HS65_LS_IVX2 U18709 ( .A(key[41]), .Z(n761) );
  HS65_LS_OAI22X1 U18710 ( .A(n768), .B(n9862), .C(n1078), .D(ld), .Z(w2[2])
         );
  HS65_LS_IVX2 U18711 ( .A(key[34]), .Z(n768) );
  HS65_LS_OAI22X1 U18712 ( .A(n764), .B(n9862), .C(n1070), .D(ld), .Z(w2[6])
         );
  HS65_LS_IVX2 U18713 ( .A(key[38]), .Z(n764) );
  HS65_LS_OAI22X1 U18714 ( .A(n759), .B(n9862), .C(n1060), .D(n9854), .Z(
        w2[11]) );
  HS65_LS_IVX2 U18715 ( .A(key[43]), .Z(n759) );
  HS65_LS_OAI22X1 U18716 ( .A(n766), .B(n9862), .C(n1074), .D(n9847), .Z(w2[4]) );
  HS65_LS_IVX2 U18717 ( .A(key[36]), .Z(n766) );
  HS65_LS_OAI22X1 U18718 ( .A(n758), .B(n9862), .C(n1058), .D(n9846), .Z(
        w2[12]) );
  HS65_LS_IVX2 U18719 ( .A(key[44]), .Z(n758) );
  HS65_LS_OAI22X1 U18720 ( .A(n765), .B(n9862), .C(n1072), .D(n9848), .Z(w2[5]) );
  HS65_LS_IVX2 U18721 ( .A(key[37]), .Z(n765) );
  HS65_LS_OAI22X1 U18722 ( .A(n757), .B(n9862), .C(n1056), .D(n9846), .Z(
        w2[13]) );
  HS65_LS_IVX2 U18723 ( .A(key[45]), .Z(n757) );
  HS65_LS_OAI22X1 U18724 ( .A(n769), .B(n9862), .C(n1080), .D(n9850), .Z(w2[1]) );
  HS65_LS_IVX2 U18725 ( .A(key[33]), .Z(n769) );
  HS65_LS_OAI22X1 U18726 ( .A(n756), .B(n9862), .C(n1054), .D(ld), .Z(w2[14])
         );
  HS65_LS_IVX2 U18727 ( .A(key[46]), .Z(n756) );
  HS65_LS_OAI22X1 U18728 ( .A(n739), .B(n9866), .C(n1020), .D(ld), .Z(w2[31])
         );
  HS65_LS_IVX2 U18729 ( .A(key[63]), .Z(n739) );
  HS65_LS_OAI22X1 U18730 ( .A(n770), .B(n9861), .C(n1082), .D(n9846), .Z(w2[0]) );
  HS65_LS_IVX2 U18731 ( .A(key[32]), .Z(n770) );
  HS65_LS_OAI22X1 U18732 ( .A(n746), .B(n9861), .C(n1034), .D(ld), .Z(w2[24])
         );
  HS65_LS_IVX2 U18733 ( .A(key[56]), .Z(n746) );
  HS65_LS_OAI22X1 U18734 ( .A(n747), .B(n9865), .C(n1036), .D(n9846), .Z(
        w2[23]) );
  HS65_LS_IVX2 U18735 ( .A(key[55]), .Z(n747) );
  HS65_LS_OAI22X1 U18736 ( .A(n745), .B(n9861), .C(n1032), .D(n9851), .Z(
        w2[25]) );
  HS65_LS_IVX2 U18737 ( .A(key[57]), .Z(n745) );
  HS65_LS_OAI22X1 U18738 ( .A(n743), .B(n9862), .C(n1028), .D(n9846), .Z(
        w2[27]) );
  HS65_LS_IVX2 U18739 ( .A(key[59]), .Z(n743) );
  HS65_LS_OAI22X1 U18740 ( .A(n744), .B(n9862), .C(n1030), .D(n9846), .Z(
        w2[26]) );
  HS65_LS_IVX2 U18741 ( .A(key[58]), .Z(n744) );
  HS65_LS_OAI22X1 U18742 ( .A(n742), .B(n9861), .C(n1026), .D(n9850), .Z(
        w2[28]) );
  HS65_LS_IVX2 U18743 ( .A(key[60]), .Z(n742) );
  HS65_LS_OAI22X1 U18744 ( .A(n741), .B(n9861), .C(n1024), .D(n9846), .Z(
        w2[29]) );
  HS65_LS_IVX2 U18745 ( .A(key[61]), .Z(n741) );
  HS65_LS_OAI22X1 U18746 ( .A(n740), .B(n9865), .C(n1022), .D(ld), .Z(w2[30])
         );
  HS65_LS_IVX2 U18747 ( .A(key[62]), .Z(n740) );
  HS65_LS_OAI22X1 U18748 ( .A(n730), .B(n9862), .C(n1004), .D(n9848), .Z(
        w0[14]) );
  HS65_LS_IVX2 U18749 ( .A(key[110]), .Z(n730) );
  HS65_LS_OAI22X1 U18750 ( .A(n737), .B(n9862), .C(n1017), .D(n9850), .Z(w0[1]) );
  HS65_LS_IVX2 U18751 ( .A(key[97]), .Z(n737) );
  HS65_LS_OAI22X1 U18752 ( .A(n725), .B(n9861), .C(n996), .D(n9847), .Z(w0[22]) );
  HS65_LS_IVX2 U18753 ( .A(key[118]), .Z(n725) );
  HS65_LS_OAI22X1 U18754 ( .A(n726), .B(n9860), .C(n999), .D(n9854), .Z(w0[19]) );
  HS65_LS_IVX2 U18755 ( .A(key[115]), .Z(n726) );
  HS65_LS_OAI22X1 U18756 ( .A(n731), .B(n9861), .C(n1007), .D(n9851), .Z(
        w0[11]) );
  HS65_LS_IVX2 U18757 ( .A(key[107]), .Z(n731) );
  HS65_LS_OAI22X1 U18758 ( .A(n735), .B(n9861), .C(n1012), .D(n9848), .Z(w0[6]) );
  HS65_LS_IVX2 U18759 ( .A(key[102]), .Z(n735) );
  HS65_LS_OAI22X1 U18760 ( .A(n727), .B(n9860), .C(n1001), .D(n9850), .Z(
        w0[17]) );
  HS65_LS_IVX2 U18761 ( .A(key[113]), .Z(n727) );
  HS65_LS_OAI22X1 U18762 ( .A(n729), .B(n9860), .C(n1003), .D(ld), .Z(w0[15])
         );
  HS65_LS_IVX2 U18763 ( .A(key[111]), .Z(n729) );
  HS65_LS_OAI22X1 U18764 ( .A(n721), .B(n9859), .C(n991), .D(n9847), .Z(w0[27]) );
  HS65_LS_IVX2 U18765 ( .A(key[123]), .Z(n721) );
  HS65_LS_OAI22X1 U18766 ( .A(n732), .B(n9866), .C(n1009), .D(n9848), .Z(w0[9]) );
  HS65_LS_IVX2 U18767 ( .A(key[105]), .Z(n732) );
  HS65_LS_OAI22X1 U18768 ( .A(n734), .B(n9861), .C(n1011), .D(n9852), .Z(w0[7]) );
  HS65_LS_IVX2 U18769 ( .A(key[103]), .Z(n734) );
  HS65_LS_OAI22X1 U18770 ( .A(n722), .B(n9859), .C(n993), .D(n9847), .Z(w0[25]) );
  HS65_LS_IVX2 U18771 ( .A(key[121]), .Z(n722) );
  HS65_LS_OAI22X1 U18772 ( .A(n724), .B(n9861), .C(n995), .D(n9852), .Z(w0[23]) );
  HS65_LS_IVX2 U18773 ( .A(key[119]), .Z(n724) );
  HS65_LS_OAI22X1 U18774 ( .A(n723), .B(n9861), .C(n994), .D(n9854), .Z(w0[24]) );
  HS65_LS_IVX2 U18775 ( .A(key[120]), .Z(n723) );
  HS65_LS_OAI22X1 U18776 ( .A(n728), .B(n9859), .C(n1002), .D(n9847), .Z(
        w0[16]) );
  HS65_LS_IVX2 U18777 ( .A(key[112]), .Z(n728) );
  HS65_LS_OAI22X1 U18778 ( .A(n733), .B(n9865), .C(n1010), .D(n9852), .Z(w0[8]) );
  HS65_LS_IVX2 U18779 ( .A(key[104]), .Z(n733) );
  HS65_LS_OAI22X1 U18780 ( .A(n738), .B(n9862), .C(n1018), .D(n9851), .Z(w0[0]) );
  HS65_LS_IVX2 U18781 ( .A(key[96]), .Z(n738) );
  HS65_LS_OAI22X1 U18782 ( .A(n754), .B(n9861), .C(n1050), .D(ld), .Z(w2[16])
         );
  HS65_LS_IVX2 U18783 ( .A(key[48]), .Z(n754) );
  HS65_LS_OAI22X1 U18784 ( .A(n752), .B(n9862), .C(n1046), .D(n9846), .Z(
        w2[18]) );
  HS65_LS_IVX2 U18785 ( .A(key[50]), .Z(n752) );
  HS65_LS_OAI22X1 U18786 ( .A(n755), .B(n9861), .C(n1052), .D(n9851), .Z(
        w2[15]) );
  HS65_LS_IVX2 U18787 ( .A(key[47]), .Z(n755) );
  HS65_LS_OAI22X1 U18788 ( .A(n753), .B(n9860), .C(n1048), .D(n9846), .Z(
        w2[17]) );
  HS65_LS_IVX2 U18789 ( .A(key[49]), .Z(n753) );
  HS65_LS_OAI22X1 U18790 ( .A(n751), .B(n9860), .C(n1044), .D(ld), .Z(w2[19])
         );
  HS65_LS_IVX2 U18791 ( .A(key[51]), .Z(n751) );
  HS65_LS_OAI22X1 U18792 ( .A(n750), .B(n9865), .C(n1042), .D(n9846), .Z(
        w2[20]) );
  HS65_LS_IVX2 U18793 ( .A(key[52]), .Z(n750) );
  HS65_LS_OAI22X1 U18794 ( .A(n748), .B(n9859), .C(n1038), .D(ld), .Z(w2[22])
         );
  HS65_LS_IVX2 U18795 ( .A(key[54]), .Z(n748) );
  HS65_LS_OAI22X1 U18796 ( .A(n749), .B(n9866), .C(n1040), .D(n9847), .Z(
        w2[21]) );
  HS65_LS_IVX2 U18797 ( .A(key[53]), .Z(n749) );
  HS65_LSS_XOR2X3 U18798 ( .A(n2780), .B(n953), .Z(n9746) );
  HS65_LS_OAI22X1 U18799 ( .A(n9859), .B(n719), .C(n987), .D(n9847), .Z(w0[31]) );
  HS65_LS_IVX2 U18800 ( .A(key[127]), .Z(n719) );
  HS65_LSS_XOR3X2 U18801 ( .A(n970), .B(n9410), .C(n1115), .Z(n987) );
  HS65_LS_NAND4ABX3 U18802 ( .A(n1116), .B(n1117), .C(n1118), .D(n1119), .Z(
        n1115) );
  HS65_LS_NAND4ABX3 U18803 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .Z(
        n1116) );
  HS65_LS_OAI212X3 U18804 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .E(
        n1131), .Z(n1117) );
  HS65_LSS_XOR3X2 U18805 ( .A(n963), .B(n9163), .C(n1431), .Z(n994) );
  HS65_LS_NAND4ABX3 U18806 ( .A(n1432), .B(n1433), .C(n1434), .D(n1435), .Z(
        n1431) );
  HS65_LS_MX41X4 U18807 ( .D0(n866), .S0(n883), .D1(n867), .S1(n875), .D2(n886), .S2(n859), .D3(n887), .S3(n1178), .Z(n1433) );
  HS65_LS_NOR4ABX2 U18808 ( .A(n1176), .B(n1311), .C(n1436), .D(n1325), .Z(
        n1435) );
  HS65_LSS_XOR3X2 U18809 ( .A(n969), .B(n9425), .C(n1142), .Z(n988) );
  HS65_LS_NAND4ABX3 U18810 ( .A(n1143), .B(n1144), .C(n1145), .D(n1146), .Z(
        n1142) );
  HS65_LS_CBI4I1X3 U18811 ( .A(n1158), .B(n1128), .C(n1159), .D(n1160), .Z(
        n1143) );
  HS65_LS_AOI212X2 U18812 ( .A(n887), .B(n853), .C(n884), .D(n865), .E(n1152), 
        .Z(n1145) );
  HS65_LSS_XOR2X3 U18813 ( .A(n2808), .B(n9266), .Z(n9734) );
  HS65_LSS_XOR2X3 U18814 ( .A(n3010), .B(n9277), .Z(n9787) );
  HS65_LSS_XOR2X3 U18815 ( .A(n2768), .B(n9294), .Z(n9806) );
  HS65_LSS_XOR2X3 U18816 ( .A(n2812), .B(n9252), .Z(n9794) );
  HS65_LSS_XOR2X3 U18817 ( .A(n3011), .B(n9278), .Z(n9786) );
  HS65_LSS_XOR2X3 U18818 ( .A(n3014), .B(n9274), .Z(n9783) );
  HS65_LSS_XOR2X3 U18819 ( .A(n3543), .B(n9331), .Z(n9719) );
  HS65_LSS_XOR2X3 U18820 ( .A(n2826), .B(n9267), .Z(n9732) );
  HS65_LSS_XOR2X3 U18821 ( .A(n2822), .B(n9202), .Z(n9760) );
  HS65_LSS_XOR2X3 U18822 ( .A(n2778), .B(n9272), .Z(n9748) );
  HS65_LSS_XOR2X3 U18823 ( .A(n2810), .B(n9253), .Z(n9796) );
  HS65_LSS_XOR2X3 U18824 ( .A(n2809), .B(n9256), .Z(n9797) );
  HS65_LSS_XOR2X3 U18825 ( .A(n2830), .B(n9199), .Z(n9728) );
  HS65_LSS_XOR2X3 U18826 ( .A(n2825), .B(n9259), .Z(n9733) );
  HS65_LSS_XOR3X2 U18827 ( .A(n1202), .B(n9405), .C(n967), .Z(n990) );
  HS65_LS_NOR3X1 U18828 ( .A(n1203), .B(n1204), .C(n1205), .Z(n1202) );
  HS65_LS_OAI212X3 U18829 ( .A(n1206), .B(n1130), .C(n1207), .D(n1208), .E(
        n1209), .Z(n1205) );
  HS65_LS_NAND4ABX3 U18830 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .Z(
        n1204) );
  HS65_LSS_XOR3X2 U18831 ( .A(n1161), .B(n9165), .C(n968), .Z(n989) );
  HS65_LS_NOR3X1 U18832 ( .A(n1162), .B(n1163), .C(n1164), .Z(n1161) );
  HS65_LS_NAND4ABX3 U18833 ( .A(n1189), .B(n1190), .C(n1191), .D(n1192), .Z(
        n1162) );
  HS65_LS_OAI212X3 U18834 ( .A(n1129), .B(n1134), .C(n1156), .D(n1186), .E(
        n1187), .Z(n1163) );
  HS65_LSS_XOR3X2 U18835 ( .A(n966), .B(n9162), .C(n1265), .Z(n991) );
  HS65_LS_NAND4ABX3 U18836 ( .A(n1266), .B(n1267), .C(n1268), .D(n1269), .Z(
        n1265) );
  HS65_LS_MX41X4 U18837 ( .D0(n856), .S0(n880), .D1(n884), .S1(n868), .D2(n854), .S2(n875), .D3(n886), .S3(n1178), .Z(n1267) );
  HS65_LS_AOI212X2 U18838 ( .A(n869), .B(n1270), .C(n885), .D(n1247), .E(n1271), .Z(n1269) );
  HS65_LSS_XOR3X2 U18839 ( .A(n964), .B(n9406), .C(n1406), .Z(n993) );
  HS65_LS_NAND4ABX3 U18840 ( .A(n1407), .B(n1408), .C(n1409), .D(n1410), .Z(
        n1406) );
  HS65_LS_AOI222X2 U18841 ( .A(n877), .B(n855), .C(n874), .D(n1429), .E(n886), 
        .F(n854), .Z(n1409) );
  HS65_LS_CB4I6X4 U18842 ( .A(n858), .B(n863), .C(n885), .D(n1327), .Z(n1407)
         );
  HS65_LSS_XOR3X2 U18843 ( .A(n2645), .B(n9170), .C(n2646), .Z(n2643) );
  HS65_LSS_XOR3X2 U18844 ( .A(n2770), .B(n9204), .C(n2817), .Z(n5976) );
  HS65_LSS_XOR3X2 U18845 ( .A(n2823), .B(n9205), .C(n275), .Z(n5949) );
  HS65_LS_OAI22X1 U18846 ( .A(n2708), .B(n9144), .C(n9141), .D(n2709), .Z(
        sa13[3]) );
  HS65_LSS_XOR2X3 U18847 ( .A(n873), .B(n9608), .Z(n2708) );
  HS65_LSS_XOR3X2 U18848 ( .A(n2704), .B(n2710), .C(n2711), .Z(n2709) );
  HS65_LSS_XOR3X2 U18849 ( .A(n873), .B(n2673), .C(n2712), .Z(n2710) );
  HS65_LS_OAI22X1 U18850 ( .A(n4421), .B(n9148), .C(n9139), .D(n4422), .Z(
        sa20[7]) );
  HS65_LSS_XOR2X3 U18851 ( .A(n957), .B(n9700), .Z(n4421) );
  HS65_LSS_XOR3X2 U18852 ( .A(n2807), .B(n4423), .C(n4424), .Z(n4422) );
  HS65_LSS_XOR3X2 U18853 ( .A(n2783), .B(n957), .C(n2784), .Z(n4423) );
  HS65_LS_OAI22X1 U18854 ( .A(n2702), .B(n9144), .C(n9141), .D(n2703), .Z(
        sa13[4]) );
  HS65_LSS_XOR2X3 U18855 ( .A(n890), .B(n9609), .Z(n2702) );
  HS65_LSS_XOR3X2 U18856 ( .A(n2704), .B(n2705), .C(n2706), .Z(n2703) );
  HS65_LSS_XOR3X2 U18857 ( .A(n890), .B(n2666), .C(n2707), .Z(n2705) );
  HS65_LS_OAI22X1 U18858 ( .A(n4810), .B(n9144), .C(n9138), .D(n4811), .Z(
        sa30[4]) );
  HS65_LSS_XOR2X3 U18859 ( .A(n954), .B(n9689), .Z(n4810) );
  HS65_LSS_XOR3X2 U18860 ( .A(n4408), .B(n4812), .C(n4813), .Z(n4811) );
  HS65_LSS_XOR3X2 U18861 ( .A(n954), .B(n4369), .C(n3224), .Z(n4812) );
  HS65_LS_OAI22X1 U18862 ( .A(n9437), .B(n9580), .C(n9587), .D(n9414), .Z(
        sa33[3]) );
  HS65_LSS_XOR2X3 U18863 ( .A(n791), .B(n9592), .Z(n3545) );
  HS65_LSS_XOR3X2 U18864 ( .A(n2715), .B(n3547), .C(n3229), .Z(n3546) );
  HS65_LSS_XOR3X2 U18865 ( .A(n791), .B(n2666), .C(n2659), .Z(n3547) );
  HS65_LS_OAI22X1 U18866 ( .A(n7562), .B(n9142), .C(n9139), .D(n7563), .Z(
        sa02[2]) );
  HS65_LSS_XOR2X3 U18867 ( .A(n941), .B(n9647), .Z(n7562) );
  HS65_LSS_XOR3X2 U18868 ( .A(n362), .B(n7564), .C(n7565), .Z(n7563) );
  HS65_LSS_XOR3X2 U18869 ( .A(n2630), .B(n941), .C(n2810), .Z(n7564) );
  HS65_LS_OAI22X1 U18870 ( .A(n5571), .B(n9143), .C(n9138), .D(n5572), .Z(
        sa30[1]) );
  HS65_LSS_XOR2X3 U18871 ( .A(n952), .B(n9686), .Z(n5571) );
  HS65_LSS_XOR3X2 U18872 ( .A(n4419), .B(n5573), .C(n4813), .Z(n5572) );
  HS65_LSS_XOR3X2 U18873 ( .A(n952), .B(n4382), .C(n3221), .Z(n5573) );
  HS65_LS_OAI22X1 U18874 ( .A(n2718), .B(n9144), .C(n9141), .D(n2719), .Z(
        sa13[1]) );
  HS65_LSS_XOR2X3 U18875 ( .A(n871), .B(n9606), .Z(n2718) );
  HS65_LSS_XOR3X2 U18876 ( .A(n2704), .B(n2720), .C(n2721), .Z(n2719) );
  HS65_LSS_XOR3X2 U18877 ( .A(n871), .B(n2685), .C(n2722), .Z(n2720) );
  HS65_LSS_XOR3X2 U18878 ( .A(n9264), .B(n2777), .C(n2801), .Z(n4445) );
  HS65_LSS_XOR3X2 U18879 ( .A(n9221), .B(n2769), .C(n2793), .Z(n6038) );
  HS65_LS_OAI22X1 U18880 ( .A(n7589), .B(n9142), .C(n9588), .D(n7590), .Z(
        sa12[3]) );
  HS65_LSS_XOR2X3 U18881 ( .A(n939), .B(n9640), .Z(n7589) );
  HS65_LSS_XOR3X2 U18882 ( .A(n7586), .B(n7591), .C(n7592), .Z(n7590) );
  HS65_LSS_XOR3X2 U18883 ( .A(n939), .B(n7565), .C(n2788), .Z(n7591) );
  HS65_LS_OAI22X1 U18884 ( .A(n7597), .B(n9142), .C(n9139), .D(n7598), .Z(
        sa12[1]) );
  HS65_LSS_XOR2X3 U18885 ( .A(n937), .B(n9638), .Z(n7597) );
  HS65_LSS_XOR3X2 U18886 ( .A(n7586), .B(n7599), .C(n7600), .Z(n7598) );
  HS65_LSS_XOR3X2 U18887 ( .A(n937), .B(n2633), .C(n2786), .Z(n7599) );
  HS65_LS_OAI22X1 U18888 ( .A(n4413), .B(n9148), .C(n9139), .D(n4414), .Z(
        sa10[1]) );
  HS65_LSS_XOR2X3 U18889 ( .A(n959), .B(n9702), .Z(n4413) );
  HS65_LSS_XOR3X2 U18890 ( .A(n4402), .B(n4415), .C(n4416), .Z(n4414) );
  HS65_LSS_XOR3X2 U18891 ( .A(n959), .B(n4387), .C(n2802), .Z(n4415) );
  HS65_LS_OAI22X1 U18892 ( .A(n5129), .B(n9146), .C(n9138), .D(n5130), .Z(
        sa30[3]) );
  HS65_LSS_XOR2X3 U18893 ( .A(n953), .B(n9688), .Z(n5129) );
  HS65_LSS_XNOR3X2 U18894 ( .A(n4411), .B(n5131), .C(n4813), .Z(n5130) );
  HS65_LSS_XOR3X2 U18895 ( .A(n953), .B(n4374), .C(n3223), .Z(n5131) );
  HS65_LS_OAI22X1 U18896 ( .A(n9436), .B(n9578), .C(n9585), .D(n9413), .Z(
        sa32[7]) );
  HS65_LSS_XOR2X3 U18897 ( .A(n935), .B(n9628), .Z(n7785) );
  HS65_LSS_XOR3X2 U18898 ( .A(n7556), .B(n7578), .C(n7787), .Z(n7786) );
  HS65_LSS_XOR2X3 U18899 ( .A(n935), .B(n2792), .Z(n7787) );
  HS65_LS_OAI22X1 U18900 ( .A(n9435), .B(n9582), .C(n9586), .D(n9412), .Z(
        sa22[6]) );
  HS65_LSS_XNOR2X3 U18901 ( .A(n9284), .B(n9635), .Z(n7607) );
  HS65_LSS_XOR3X2 U18902 ( .A(n2815), .B(n7578), .C(n7609), .Z(n7608) );
  HS65_LSS_XOR3X2 U18903 ( .A(n2766), .B(n9284), .C(n579), .Z(n7609) );
  HS65_LS_OAI22X1 U18904 ( .A(n4358), .B(n9143), .C(n9588), .D(n4359), .Z(
        sa00[6]) );
  HS65_LSS_XOR2X3 U18905 ( .A(n969), .B(n9715), .Z(n4358) );
  HS65_LSS_XNOR3X2 U18906 ( .A(n3225), .B(n4360), .C(n4361), .Z(n4359) );
  HS65_LSS_XOR3X2 U18907 ( .A(n2783), .B(n969), .C(n2830), .Z(n4360) );
  HS65_LS_OAI22X1 U18908 ( .A(n5951), .B(n9147), .C(n9138), .D(n5952), .Z(
        sa01[6]) );
  HS65_LSS_XOR2X3 U18909 ( .A(n950), .B(n9683), .Z(n5951) );
  HS65_LSS_XNOR3X2 U18910 ( .A(n3217), .B(n5953), .C(n5954), .Z(n5952) );
  HS65_LSS_XOR3X2 U18911 ( .A(n2775), .B(n950), .C(n2822), .Z(n5953) );
  HS65_LS_OAI22X1 U18912 ( .A(n9434), .B(n9582), .C(n9584), .D(n9411), .Z(
        sa02[6]) );
  HS65_LSS_XOR2X3 U18913 ( .A(n943), .B(n9651), .Z(n7543) );
  HS65_LSS_XOR3X2 U18914 ( .A(n3013), .B(n7545), .C(n7546), .Z(n7544) );
  HS65_LSS_XOR3X2 U18915 ( .A(n2767), .B(n943), .C(n2814), .Z(n7546) );
  HS65_LS_AO22X4 U18916 ( .A(key[88]), .B(n9857), .C(n1090), .D(n9860), .Z(
        w1[24]) );
  HS65_LS_AO22X4 U18917 ( .A(key[86]), .B(n9858), .C(n1092), .D(n9864), .Z(
        w1[22]) );
  HS65_LS_AO22X4 U18918 ( .A(key[72]), .B(n9855), .C(n1106), .D(n9866), .Z(
        w1[8]) );
  HS65_LS_AO22X4 U18919 ( .A(key[87]), .B(n9857), .C(n1091), .D(n9864), .Z(
        w1[23]) );
  HS65_LS_AO22X4 U18920 ( .A(key[80]), .B(n9854), .C(n1098), .D(n9866), .Z(
        w1[16]) );
  HS65_LS_AO22X4 U18921 ( .A(key[71]), .B(n9858), .C(n1107), .D(n9866), .Z(
        w1[7]) );
  HS65_LS_AO22X4 U18922 ( .A(key[64]), .B(n9857), .C(n1114), .D(n9866), .Z(
        w1[0]) );
  HS65_LS_AO22X4 U18923 ( .A(key[70]), .B(n9855), .C(n1108), .D(n9863), .Z(
        w1[6]) );
  HS65_LS_AO22X4 U18924 ( .A(key[101]), .B(n9856), .C(n1013), .D(n9864), .Z(
        w0[5]) );
  HS65_LS_AO22X4 U18925 ( .A(key[98]), .B(n9856), .C(n1016), .D(n9864), .Z(
        w0[2]) );
  HS65_LS_AO22X4 U18926 ( .A(key[78]), .B(n9858), .C(n1100), .D(n9866), .Z(
        w1[14]) );
  HS65_LS_AO22X4 U18927 ( .A(key[65]), .B(n9854), .C(n1113), .D(n9859), .Z(
        w1[1]) );
  HS65_LS_AO22X4 U18928 ( .A(key[67]), .B(n9855), .C(n1111), .D(n9865), .Z(
        w1[3]) );
  HS65_LS_AO22X4 U18929 ( .A(key[73]), .B(n9858), .C(n1105), .D(n9866), .Z(
        w1[9]) );
  HS65_LS_AO22X4 U18930 ( .A(key[91]), .B(n9857), .C(n1087), .D(n9863), .Z(
        w1[27]) );
  HS65_LS_AO22X4 U18931 ( .A(key[81]), .B(n9854), .C(n1097), .D(n9866), .Z(
        w1[17]) );
  HS65_LS_AO22X4 U18932 ( .A(key[83]), .B(n9855), .C(n1095), .D(n9866), .Z(
        w1[19]) );
  HS65_LS_AO22X4 U18933 ( .A(key[79]), .B(n9858), .C(n1099), .D(n9866), .Z(
        w1[15]) );
  HS65_LS_AO22X4 U18934 ( .A(key[75]), .B(n9855), .C(n1103), .D(n9866), .Z(
        w1[11]) );
  HS65_LS_AO22X4 U18935 ( .A(key[109]), .B(n9855), .C(n1005), .D(n9866), .Z(
        w0[13]) );
  HS65_LS_AO22X4 U18936 ( .A(key[108]), .B(n9855), .C(n1006), .D(n9864), .Z(
        w0[12]) );
  HS65_LS_AO22X4 U18937 ( .A(key[66]), .B(n9854), .C(n1112), .D(n9859), .Z(
        w1[2]) );
  HS65_LS_AO22X4 U18938 ( .A(key[69]), .B(n9858), .C(n1109), .D(n9859), .Z(
        w1[5]) );
  HS65_LS_AO22X4 U18939 ( .A(key[116]), .B(n9858), .C(n998), .D(n9864), .Z(
        w0[20]) );
  HS65_LS_AO22X4 U18940 ( .A(key[74]), .B(n9854), .C(n1104), .D(n9864), .Z(
        w1[10]) );
  HS65_LS_AO22X4 U18941 ( .A(key[77]), .B(n9854), .C(n1101), .D(n9864), .Z(
        w1[13]) );
  HS65_LS_AO22X4 U18942 ( .A(key[76]), .B(n9858), .C(n1102), .D(n9864), .Z(
        w1[12]) );
  HS65_LS_AO22X4 U18943 ( .A(key[68]), .B(n9854), .C(n1110), .D(n9859), .Z(
        w1[4]) );
  HS65_LS_AO22X4 U18944 ( .A(key[84]), .B(n9858), .C(n1094), .D(n9864), .Z(
        w1[20]) );
  HS65_LS_AO22X4 U18945 ( .A(key[95]), .B(n9857), .C(n1083), .D(n9861), .Z(
        w1[31]) );
  HS65_LS_AO22X4 U18946 ( .A(key[89]), .B(n9857), .C(n1089), .D(n9865), .Z(
        w1[25]) );
  HS65_LS_AO22X4 U18947 ( .A(key[94]), .B(n9857), .C(n1084), .D(n9865), .Z(
        w1[30]) );
  HS65_LS_AO22X4 U18948 ( .A(key[85]), .B(n9858), .C(n1093), .D(n9864), .Z(
        w1[21]) );
  HS65_LS_AO22X4 U18949 ( .A(key[100]), .B(n9856), .C(n1014), .D(n9864), .Z(
        \u0/N46 ) );
  HS65_LS_AO22X4 U18950 ( .A(key[82]), .B(n9858), .C(n1096), .D(n9864), .Z(
        w1[18]) );
  HS65_LS_AO22X4 U18951 ( .A(key[93]), .B(n9857), .C(n1085), .D(n9865), .Z(
        w1[29]) );
  HS65_LS_AO22X4 U18952 ( .A(key[117]), .B(n9857), .C(n997), .D(n9864), .Z(
        w0[21]) );
  HS65_LS_AO22X4 U18953 ( .A(key[90]), .B(n9856), .C(n1088), .D(n9865), .Z(
        w1[26]) );
  HS65_LS_AO22X4 U18954 ( .A(key[92]), .B(n9857), .C(n1086), .D(n9865), .Z(
        w1[28]) );
  HS65_LS_AO22X4 U18955 ( .A(key[106]), .B(n9858), .C(n1008), .D(n9864), .Z(
        w0[10]) );
  HS65_LS_AO22X4 U18956 ( .A(key[114]), .B(n9855), .C(n1000), .D(n9864), .Z(
        w0[18]) );
  HS65_LS_AO22X4 U18957 ( .A(key[125]), .B(n9855), .C(n989), .D(n9865), .Z(
        w0[29]) );
  HS65_LS_AO22X4 U18958 ( .A(key[124]), .B(n9855), .C(n990), .D(n9865), .Z(
        w0[28]) );
  HS65_LS_AO22X4 U18959 ( .A(key[122]), .B(n9855), .C(n992), .D(n9864), .Z(
        w0[26]) );
  HS65_LS_AO22X4 U18960 ( .A(key[0]), .B(n9857), .C(n1081), .D(n9865), .Z(
        w3[0]) );
  HS65_LSS_XOR2X3 U18961 ( .A(n788), .B(n1082), .Z(n1081) );
  HS65_LS_AO22X4 U18962 ( .A(key[2]), .B(n9857), .C(n1077), .D(n9865), .Z(
        w3[2]) );
  HS65_LSS_XOR2X3 U18963 ( .A(n790), .B(n1078), .Z(n1077) );
  HS65_LS_AO22X4 U18964 ( .A(key[8]), .B(n9857), .C(n1065), .D(n9863), .Z(
        w3[8]) );
  HS65_LSS_XOR2X3 U18965 ( .A(n829), .B(n1066), .Z(n1065) );
  HS65_LS_AO22X4 U18966 ( .A(key[6]), .B(n9857), .C(n1069), .D(n9863), .Z(
        w3[6]) );
  HS65_LSS_XOR2X3 U18967 ( .A(n810), .B(n1070), .Z(n1069) );
  HS65_LS_AO22X4 U18968 ( .A(key[24]), .B(n9856), .C(n1033), .D(n9865), .Z(
        w3[24]) );
  HS65_LSS_XOR2X3 U18969 ( .A(n911), .B(n1034), .Z(n1033) );
  HS65_LS_AO22X4 U18970 ( .A(key[4]), .B(n9857), .C(n1073), .D(n9863), .Z(
        w3[4]) );
  HS65_LSS_XOR2X3 U18971 ( .A(n808), .B(n1074), .Z(n1073) );
  HS65_LS_AO22X4 U18972 ( .A(key[12]), .B(n9857), .C(n1057), .D(n9863), .Z(
        w3[12]) );
  HS65_LSS_XOR2X3 U18973 ( .A(n849), .B(n1058), .Z(n1057) );
  HS65_LS_AO22X4 U18974 ( .A(key[10]), .B(n9857), .C(n1061), .D(n9863), .Z(
        w3[10]) );
  HS65_LSS_XOR2X3 U18975 ( .A(n831), .B(n1062), .Z(n1061) );
  HS65_LS_AO22X4 U18976 ( .A(key[31]), .B(n9856), .C(n1019), .D(n9863), .Z(
        w3[31]) );
  HS65_LSS_XOR2X3 U18977 ( .A(n934), .B(n1020), .Z(n1019) );
  HS65_LS_AO22X4 U18978 ( .A(key[14]), .B(n9858), .C(n1053), .D(n9863), .Z(
        w3[14]) );
  HS65_LSS_XOR2X3 U18979 ( .A(n851), .B(n1054), .Z(n1053) );
  HS65_LS_AO22X4 U18980 ( .A(key[29]), .B(n9856), .C(n1023), .D(n9863), .Z(
        w3[29]) );
  HS65_LSS_XOR2X3 U18981 ( .A(n932), .B(n1024), .Z(n1023) );
  HS65_LS_AO22X4 U18982 ( .A(key[3]), .B(n9858), .C(n1075), .D(n9863), .Z(
        w3[3]) );
  HS65_LSS_XOR2X3 U18983 ( .A(n791), .B(n1076), .Z(n1075) );
  HS65_LS_AO22X4 U18984 ( .A(key[28]), .B(n9856), .C(n1025), .D(n9863), .Z(
        w3[28]) );
  HS65_LSS_XOR2X3 U18985 ( .A(n931), .B(n1026), .Z(n1025) );
  HS65_LS_AO22X4 U18986 ( .A(key[1]), .B(n9858), .C(n1079), .D(n9863), .Z(
        w3[1]) );
  HS65_LSS_XOR2X3 U18987 ( .A(n789), .B(n1080), .Z(n1079) );
  HS65_LS_AO22X4 U18988 ( .A(key[11]), .B(n9858), .C(n1059), .D(n9863), .Z(
        w3[11]) );
  HS65_LSS_XOR2X3 U18989 ( .A(n832), .B(n1060), .Z(n1059) );
  HS65_LS_AO22X4 U18990 ( .A(key[9]), .B(n9854), .C(n1063), .D(n9859), .Z(
        w3[9]) );
  HS65_LSS_XOR2X3 U18991 ( .A(n830), .B(n1064), .Z(n1063) );
  HS65_LS_AO22X4 U18992 ( .A(key[20]), .B(n9856), .C(n1041), .D(n9863), .Z(
        w3[20]) );
  HS65_LSS_XOR2X3 U18993 ( .A(n890), .B(n1042), .Z(n1041) );
  HS65_LS_AO22X4 U18994 ( .A(key[18]), .B(n9856), .C(n1045), .D(n9859), .Z(
        w3[18]) );
  HS65_LSS_XOR2X3 U18995 ( .A(n872), .B(n1046), .Z(n1045) );
  HS65_LS_AO22X4 U18996 ( .A(key[16]), .B(n9858), .C(n1049), .D(n9866), .Z(
        w3[16]) );
  HS65_LSS_XOR2X3 U18997 ( .A(n870), .B(n1050), .Z(n1049) );
  HS65_LS_AO22X4 U18998 ( .A(key[21]), .B(n9856), .C(n1039), .D(n9863), .Z(
        w3[21]) );
  HS65_LSS_XOR2X3 U18999 ( .A(n891), .B(n1040), .Z(n1039) );
  HS65_LS_AO22X4 U19000 ( .A(key[7]), .B(n9858), .C(n1067), .D(n9866), .Z(
        w3[7]) );
  HS65_LSS_XOR2X3 U19001 ( .A(n811), .B(n1068), .Z(n1067) );
  HS65_LS_AO22X4 U19002 ( .A(key[30]), .B(n9856), .C(n1021), .D(n9863), .Z(
        w3[30]) );
  HS65_LSS_XOR2X3 U19003 ( .A(n933), .B(n1022), .Z(n1021) );
  HS65_LS_AO22X4 U19004 ( .A(key[26]), .B(n9855), .C(n1029), .D(n9863), .Z(
        w3[26]) );
  HS65_LSS_XOR2X3 U19005 ( .A(n913), .B(n1030), .Z(n1029) );
  HS65_LS_AO22X4 U19006 ( .A(key[19]), .B(n9855), .C(n1043), .D(n9863), .Z(
        w3[19]) );
  HS65_LSS_XOR2X3 U19007 ( .A(n873), .B(n1044), .Z(n1043) );
  HS65_LS_AO22X4 U19008 ( .A(key[17]), .B(n9855), .C(n1047), .D(n9859), .Z(
        w3[17]) );
  HS65_LSS_XOR2X3 U19009 ( .A(n871), .B(n1048), .Z(n1047) );
  HS65_LS_AO22X4 U19010 ( .A(key[27]), .B(n9855), .C(n1027), .D(n9863), .Z(
        w3[27]) );
  HS65_LSS_XOR2X3 U19011 ( .A(n914), .B(n1028), .Z(n1027) );
  HS65_LSS_XOR2X3 U19012 ( .A(n9579), .B(n9577), .Z(n978) );
  HS65_LS_IVX2 U19013 ( .A(n9577), .Z(n972) );
  HS65_LS_OAI211X5 U19014 ( .A(n9164), .B(n3), .C(rst), .D(n9860), .Z(n2619)
         );
  HS65_LS_NAND2X2 U19015 ( .A(n984), .B(n9577), .Z(n983) );
  HS65_LS_OAI32X2 U19016 ( .A(n975), .B(n9577), .C(n982), .D(n9846), .E(n983), 
        .Z(\u0/rcon [27]) );
  HS65_LSS_XOR2X3 U19017 ( .A(n985), .B(n9571), .Z(n974) );
  HS65_LS_NAND2X2 U19018 ( .A(n9572), .B(n986), .Z(n985) );
  HS65_LS_IVX2 U19019 ( .A(n9259), .Z(n958) );
  HS65_LS_IVX2 U19020 ( .A(n9256), .Z(n936) );
  HS65_LS_IVX2 U19021 ( .A(n9294), .Z(n935) );
  HS65_LS_IVX2 U19022 ( .A(n9249), .Z(n940) );
  HS65_LS_IVX2 U19023 ( .A(n9199), .Z(n962) );
  HS65_LS_IVX2 U19024 ( .A(n9202), .Z(n945) );
  HS65_LS_NOR3X1 U19025 ( .A(n9161), .B(n9407), .C(n9408), .Z(n2623) );
  HS65_LS_IVX2 U19026 ( .A(n9266), .Z(n957) );
  HS65_LS_IVX2 U19027 ( .A(n9277), .Z(n941) );
  HS65_LS_IVX2 U19028 ( .A(n9274), .Z(n943) );
  HS65_LS_IVX4 U19029 ( .A(n9588), .Z(n9148) );
  HS65_LS_IVX2 U19030 ( .A(n9272), .Z(n952) );
  HS65_LS_IVX2 U19031 ( .A(n9267), .Z(n959) );
  HS65_LS_IVX2 U19032 ( .A(n9278), .Z(n942) );
  HS65_LS_IVX2 U19033 ( .A(n9253), .Z(n937) );
  HS65_LS_IVX2 U19034 ( .A(n9252), .Z(n939) );
  HS65_LS_IVX2 U19035 ( .A(n9255), .Z(n938) );
  HS65_LSS_XNOR2X3 U19036 ( .A(n986), .B(n9572), .Z(n981) );
  HS65_LS_OAI13X1 U19037 ( .A(n978), .B(n9577), .C(n977), .D(n979), .Z(
        \u0/rcon [29]) );
  HS65_LS_IVX2 U19038 ( .A(n9195), .Z(n960) );
  HS65_LS_IVX2 U19039 ( .A(n9273), .Z(n956) );
  HS65_LS_IVX2 U19040 ( .A(n9201), .Z(n944) );
  HS65_LS_IVX2 U19041 ( .A(n9331), .Z(n969) );
  HS65_LS_IVX2 U19042 ( .A(n9270), .Z(n961) );
  HS65_LS_IVX2 U19043 ( .A(n9196), .Z(n955) );
  HS65_LS_IVX2 U19044 ( .A(n9198), .Z(n947) );
  HS65_LS_IVX2 U19045 ( .A(n9200), .Z(n949) );
  HS65_LSS_XOR2X3 U19046 ( .A(n9289), .B(n2765), .Z(n9809) );
  HS65_LS_IVX2 U19047 ( .A(n9197), .Z(n948) );
  HS65_LS_IVX2 U19048 ( .A(n9203), .Z(n950) );
  HS65_LS_IVX2 U19049 ( .A(n9260), .Z(n963) );
  HS65_LSS_XOR2X3 U19050 ( .A(n2790), .B(n9286), .Z(n9800) );
  HS65_LSS_XOR2X3 U19051 ( .A(n2789), .B(n9288), .Z(n9801) );
  HS65_LS_IVX2 U19052 ( .A(n9248), .Z(n970) );
  HS65_LS_IVX2 U19053 ( .A(n9262), .Z(n964) );
  HS65_LS_IVX2 U19054 ( .A(n9265), .Z(n966) );
  HS65_LS_NOR3X1 U19055 ( .A(n977), .B(n9577), .C(n971), .Z(\u0/rcon [31]) );
  HS65_LS_IVX2 U19056 ( .A(n9192), .Z(n965) );
  HS65_LS_IVX2 U19057 ( .A(n9194), .Z(n968) );
  HS65_LS_IVX2 U19058 ( .A(n9193), .Z(n967) );
  HS65_LS_IVX2 U19059 ( .A(n9408), .Z(n5) );
  HS65_LSS_XOR2X3 U19060 ( .A(n2740), .B(n9186), .Z(n9841) );
  HS65_LSS_XOR2X3 U19061 ( .A(n2745), .B(n9175), .Z(n9825) );
  HS65_LSS_XOR2X3 U19062 ( .A(n2652), .B(n9393), .Z(n9840) );
  HS65_LSS_XOR2X3 U19063 ( .A(n2647), .B(n9172), .Z(n9824) );
  HS65_LS_OAI31X5 U19064 ( .A(n1), .B(n2623), .C(n2619), .D(n2622), .Z(dcnt[3]) );
  HS65_LS_IVX2 U19065 ( .A(n9164), .Z(n1) );
  HS65_LS_NAND2X7 U19066 ( .A(n9846), .B(rst), .Z(n2622) );
  HS65_LS_NOR3AX2 U19067 ( .A(n9135), .B(n9161), .C(n5), .Z(n9717) );
  HS65_LS_NOR3X1 U19068 ( .A(n9407), .B(n9164), .C(n9847), .Z(n9135) );
  HS65_LSS_XOR2X3 U19069 ( .A(n2814), .B(n9249), .Z(n9792) );
  HS65_LS_OAI21X3 U19070 ( .A(n9408), .B(n2619), .C(n2622), .Z(dcnt[0]) );
  HS65_LS_OAI21X3 U19071 ( .A(n3), .B(n2619), .C(n2620), .Z(dcnt[2]) );
  HS65_LS_CBI4I1X5 U19072 ( .A(n9161), .B(n2), .C(n2621), .D(n9407), .Z(n2620)
         );
  HS65_LS_AND2X4 U19073 ( .A(n9579), .B(n9577), .Z(n986) );
  HS65_LS_AO312X9 U19074 ( .A(n5), .B(n4), .C(n2), .D(n2621), .E(n9161), .F(
        n715), .Z(dcnt[1]) );
  HS65_LS_IVX2 U19075 ( .A(n9161), .Z(n4) );
  HS65_LS_IVX9 U19076 ( .A(n2622), .Z(n715) );
  HS65_LS_DFPHQX4 clk_r_REG430_S1 ( .D(text_in_r[127]), .E(n9847), .CP(clk), 
        .Q(n9716) );
  HS65_LS_DFPHQX4 clk_r_REG431_S1 ( .D(text_in_r[126]), .E(n9847), .CP(clk), 
        .Q(n9715) );
  HS65_LS_DFPHQX4 clk_r_REG432_S1 ( .D(text_in_r[125]), .E(n9847), .CP(clk), 
        .Q(n9714) );
  HS65_LS_DFPHQX4 clk_r_REG433_S1 ( .D(text_in_r[124]), .E(n9847), .CP(clk), 
        .Q(n9713) );
  HS65_LS_DFPHQX4 clk_r_REG434_S1 ( .D(text_in_r[123]), .E(n9847), .CP(clk), 
        .Q(n9712) );
  HS65_LS_DFPHQX4 clk_r_REG435_S1 ( .D(text_in_r[122]), .E(n9847), .CP(clk), 
        .Q(n9711) );
  HS65_LS_DFPHQX4 clk_r_REG436_S1 ( .D(text_in_r[121]), .E(n9847), .CP(clk), 
        .Q(n9710) );
  HS65_LS_DFPHQX4 clk_r_REG437_S1 ( .D(text_in_r[120]), .E(n9847), .CP(clk), 
        .Q(n9709) );
  HS65_LS_DFPHQX4 clk_r_REG438_S1 ( .D(text_in_r[119]), .E(n9847), .CP(clk), 
        .Q(n9708) );
  HS65_LS_DFPHQX4 clk_r_REG439_S1 ( .D(text_in_r[118]), .E(n9848), .CP(clk), 
        .Q(n9707) );
  HS65_LS_DFPHQX4 clk_r_REG440_S1 ( .D(text_in_r[117]), .E(n9848), .CP(clk), 
        .Q(n9706) );
  HS65_LS_DFPHQX4 clk_r_REG441_S1 ( .D(text_in_r[116]), .E(n9848), .CP(clk), 
        .Q(n9705) );
  HS65_LS_DFPHQX4 clk_r_REG442_S1 ( .D(text_in_r[115]), .E(n9848), .CP(clk), 
        .Q(n9704) );
  HS65_LS_DFPHQX4 clk_r_REG443_S1 ( .D(text_in_r[114]), .E(n9848), .CP(clk), 
        .Q(n9703) );
  HS65_LS_DFPHQX4 clk_r_REG444_S1 ( .D(text_in_r[113]), .E(n9848), .CP(clk), 
        .Q(n9702) );
  HS65_LS_DFPHQX4 clk_r_REG445_S1 ( .D(text_in_r[112]), .E(n9848), .CP(clk), 
        .Q(n9701) );
  HS65_LS_DFPHQX4 clk_r_REG446_S1 ( .D(text_in_r[111]), .E(n9848), .CP(clk), 
        .Q(n9700) );
  HS65_LS_DFPHQX4 clk_r_REG447_S1 ( .D(text_in_r[110]), .E(n9848), .CP(clk), 
        .Q(n9699) );
  HS65_LS_DFPHQX4 clk_r_REG448_S1 ( .D(text_in_r[109]), .E(n9848), .CP(clk), 
        .Q(n9698) );
  HS65_LS_DFPHQX4 clk_r_REG449_S1 ( .D(text_in_r[108]), .E(n9848), .CP(clk), 
        .Q(n9697) );
  HS65_LS_DFPHQX4 clk_r_REG450_S1 ( .D(text_in_r[107]), .E(n9848), .CP(clk), 
        .Q(n9696) );
  HS65_LS_DFPHQX4 clk_r_REG451_S1 ( .D(text_in_r[106]), .E(n9848), .CP(clk), 
        .Q(n9695) );
  HS65_LS_DFPHQX4 clk_r_REG452_S1 ( .D(text_in_r[105]), .E(n9848), .CP(clk), 
        .Q(n9694) );
  HS65_LS_DFPHQX4 clk_r_REG453_S1 ( .D(text_in_r[104]), .E(n9849), .CP(clk), 
        .Q(n9693) );
  HS65_LS_DFPHQX4 clk_r_REG454_S1 ( .D(text_in_r[103]), .E(n9849), .CP(clk), 
        .Q(n9692) );
  HS65_LS_DFPHQX4 clk_r_REG455_S1 ( .D(text_in_r[102]), .E(n9849), .CP(clk), 
        .Q(n9691) );
  HS65_LS_DFPHQX4 clk_r_REG456_S1 ( .D(text_in_r[101]), .E(n9849), .CP(clk), 
        .Q(n9690) );
  HS65_LS_DFPHQX4 clk_r_REG457_S1 ( .D(text_in_r[100]), .E(n9849), .CP(clk), 
        .Q(n9689) );
  HS65_LS_DFPHQX4 clk_r_REG458_S1 ( .D(text_in_r[99]), .E(n9849), .CP(clk), 
        .Q(n9688) );
  HS65_LS_DFPHQX4 clk_r_REG459_S1 ( .D(text_in_r[98]), .E(n9849), .CP(clk), 
        .Q(n9687) );
  HS65_LS_DFPHQX4 clk_r_REG460_S1 ( .D(text_in_r[97]), .E(n9849), .CP(clk), 
        .Q(n9686) );
  HS65_LS_DFPHQX4 clk_r_REG461_S1 ( .D(text_in_r[96]), .E(n9849), .CP(clk), 
        .Q(n9685) );
  HS65_LS_DFPHQX4 clk_r_REG462_S1 ( .D(text_in_r[95]), .E(n9849), .CP(clk), 
        .Q(n9684) );
  HS65_LS_DFPHQX4 clk_r_REG463_S1 ( .D(text_in_r[94]), .E(n9849), .CP(clk), 
        .Q(n9683) );
  HS65_LS_DFPHQX4 clk_r_REG464_S1 ( .D(text_in_r[93]), .E(n9849), .CP(clk), 
        .Q(n9682) );
  HS65_LS_DFPHQX4 clk_r_REG465_S1 ( .D(text_in_r[92]), .E(n9849), .CP(clk), 
        .Q(n9681) );
  HS65_LS_DFPHQX4 clk_r_REG466_S1 ( .D(text_in_r[91]), .E(n9853), .CP(clk), 
        .Q(n9680) );
  HS65_LS_DFPHQX4 clk_r_REG467_S1 ( .D(text_in_r[90]), .E(ld), .CP(clk), .Q(
        n9679) );
  HS65_LS_DFPHQX4 clk_r_REG468_S1 ( .D(text_in_r[89]), .E(n9852), .CP(clk), 
        .Q(n9678) );
  HS65_LS_DFPHQX4 clk_r_REG469_S1 ( .D(text_in_r[88]), .E(n9847), .CP(clk), 
        .Q(n9677) );
  HS65_LS_DFPHQX4 clk_r_REG470_S1 ( .D(text_in_r[87]), .E(n9846), .CP(clk), 
        .Q(n9676) );
  HS65_LS_DFPHQX4 clk_r_REG471_S1 ( .D(text_in_r[86]), .E(n9852), .CP(clk), 
        .Q(n9675) );
  HS65_LS_DFPHQX4 clk_r_REG472_S1 ( .D(text_in_r[85]), .E(n9847), .CP(clk), 
        .Q(n9674) );
  HS65_LS_DFPHQX4 clk_r_REG473_S1 ( .D(text_in_r[84]), .E(ld), .CP(clk), .Q(
        n9673) );
  HS65_LS_DFPHQX4 clk_r_REG474_S1 ( .D(text_in_r[83]), .E(n9853), .CP(clk), 
        .Q(n9672) );
  HS65_LS_DFPHQX4 clk_r_REG475_S1 ( .D(text_in_r[82]), .E(n9853), .CP(clk), 
        .Q(n9671) );
  HS65_LS_DFPHQX4 clk_r_REG476_S1 ( .D(text_in_r[81]), .E(n9850), .CP(clk), 
        .Q(n9670) );
  HS65_LS_DFPHQX4 clk_r_REG477_S1 ( .D(text_in_r[80]), .E(n9853), .CP(clk), 
        .Q(n9669) );
  HS65_LS_DFPHQX4 clk_r_REG478_S1 ( .D(text_in_r[79]), .E(n9851), .CP(clk), 
        .Q(n9668) );
  HS65_LS_DFPHQX4 clk_r_REG479_S1 ( .D(text_in_r[78]), .E(n9853), .CP(clk), 
        .Q(n9667) );
  HS65_LS_DFPHQX4 clk_r_REG480_S1 ( .D(text_in_r[77]), .E(n9848), .CP(clk), 
        .Q(n9666) );
  HS65_LS_DFPHQX4 clk_r_REG481_S1 ( .D(text_in_r[76]), .E(n9853), .CP(clk), 
        .Q(n9665) );
  HS65_LS_DFPHQX4 clk_r_REG482_S1 ( .D(text_in_r[75]), .E(n9853), .CP(clk), 
        .Q(n9664) );
  HS65_LS_DFPHQX4 clk_r_REG483_S1 ( .D(text_in_r[74]), .E(n9854), .CP(clk), 
        .Q(n9663) );
  HS65_LS_DFPHQX4 clk_r_REG484_S1 ( .D(text_in_r[73]), .E(n9849), .CP(clk), 
        .Q(n9662) );
  HS65_LS_DFPHQX4 clk_r_REG485_S1 ( .D(text_in_r[72]), .E(n9854), .CP(clk), 
        .Q(n9661) );
  HS65_LS_DFPHQX4 clk_r_REG486_S1 ( .D(text_in_r[71]), .E(n9853), .CP(clk), 
        .Q(n9660) );
  HS65_LS_DFPHQX4 clk_r_REG487_S1 ( .D(text_in_r[70]), .E(n9854), .CP(clk), 
        .Q(n9659) );
  HS65_LS_DFPHQX4 clk_r_REG488_S1 ( .D(text_in_r[69]), .E(n9853), .CP(clk), 
        .Q(n9658) );
  HS65_LS_DFPHQX4 clk_r_REG489_S1 ( .D(text_in_r[68]), .E(n9854), .CP(clk), 
        .Q(n9657) );
  HS65_LS_DFPHQX4 clk_r_REG490_S1 ( .D(text_in_r[67]), .E(n9853), .CP(clk), 
        .Q(n9656) );
  HS65_LS_DFPHQX4 clk_r_REG491_S1 ( .D(text_in_r[66]), .E(n9853), .CP(clk), 
        .Q(n9655) );
  HS65_LS_DFPHQX4 clk_r_REG492_S1 ( .D(text_in_r[65]), .E(n9853), .CP(clk), 
        .Q(n9654) );
  HS65_LS_DFPHQX4 clk_r_REG493_S1 ( .D(text_in_r[64]), .E(n9853), .CP(clk), 
        .Q(n9653) );
  HS65_LS_DFPHQX4 clk_r_REG494_S1 ( .D(text_in_r[63]), .E(n9854), .CP(clk), 
        .Q(n9652) );
  HS65_LS_DFPHQX4 clk_r_REG495_S1 ( .D(text_in_r[62]), .E(n9853), .CP(clk), 
        .Q(n9651) );
  HS65_LS_DFPHQX4 clk_r_REG496_S1 ( .D(text_in_r[61]), .E(n9853), .CP(clk), 
        .Q(n9650) );
  HS65_LS_DFPHQX4 clk_r_REG497_S1 ( .D(text_in_r[60]), .E(n9854), .CP(clk), 
        .Q(n9649) );
  HS65_LS_DFPHQX4 clk_r_REG498_S1 ( .D(text_in_r[59]), .E(n9854), .CP(clk), 
        .Q(n9648) );
  HS65_LS_DFPHQX4 clk_r_REG499_S1 ( .D(text_in_r[58]), .E(n9853), .CP(clk), 
        .Q(n9647) );
  HS65_LS_DFPHQX4 clk_r_REG500_S1 ( .D(text_in_r[57]), .E(n9853), .CP(clk), 
        .Q(n9646) );
  HS65_LS_DFPHQX4 clk_r_REG501_S1 ( .D(text_in_r[56]), .E(n9853), .CP(clk), 
        .Q(n9645) );
  HS65_LS_DFPHQX4 clk_r_REG502_S1 ( .D(text_in_r[55]), .E(n9853), .CP(clk), 
        .Q(n9644) );
  HS65_LS_DFPHQX4 clk_r_REG503_S1 ( .D(text_in_r[54]), .E(n9853), .CP(clk), 
        .Q(n9643) );
  HS65_LS_DFPHQX4 clk_r_REG504_S1 ( .D(text_in_r[53]), .E(ld), .CP(clk), .Q(
        n9642) );
  HS65_LS_DFPHQX4 clk_r_REG505_S1 ( .D(text_in_r[52]), .E(n9851), .CP(clk), 
        .Q(n9641) );
  HS65_LS_DFPHQX4 clk_r_REG506_S1 ( .D(text_in_r[51]), .E(n9849), .CP(clk), 
        .Q(n9640) );
  HS65_LS_DFPHQX4 clk_r_REG507_S1 ( .D(text_in_r[50]), .E(ld), .CP(clk), .Q(
        n9639) );
  HS65_LS_DFPHQX4 clk_r_REG508_S1 ( .D(text_in_r[49]), .E(n9850), .CP(clk), 
        .Q(n9638) );
  HS65_LS_DFPHQX4 clk_r_REG509_S1 ( .D(text_in_r[48]), .E(n9846), .CP(clk), 
        .Q(n9637) );
  HS65_LS_DFPHQX4 clk_r_REG510_S1 ( .D(text_in_r[47]), .E(ld), .CP(clk), .Q(
        n9636) );
  HS65_LS_DFPHQX4 clk_r_REG511_S1 ( .D(text_in_r[46]), .E(n9849), .CP(clk), 
        .Q(n9635) );
  HS65_LS_DFPHQX4 clk_r_REG512_S1 ( .D(text_in_r[45]), .E(ld), .CP(clk), .Q(
        n9634) );
  HS65_LS_DFPHQX4 clk_r_REG513_S1 ( .D(text_in_r[44]), .E(n9849), .CP(clk), 
        .Q(n9633) );
  HS65_LS_DFPHQX4 clk_r_REG514_S1 ( .D(text_in_r[43]), .E(n9852), .CP(clk), 
        .Q(n9632) );
  HS65_LS_DFPHQX4 clk_r_REG515_S1 ( .D(text_in_r[42]), .E(n9852), .CP(clk), 
        .Q(n9631) );
  HS65_LS_DFPHQX4 clk_r_REG516_S1 ( .D(text_in_r[41]), .E(n9852), .CP(clk), 
        .Q(n9630) );
  HS65_LS_DFPHQX4 clk_r_REG517_S1 ( .D(text_in_r[40]), .E(n9852), .CP(clk), 
        .Q(n9629) );
  HS65_LS_DFPHQX4 clk_r_REG518_S1 ( .D(text_in_r[39]), .E(n9852), .CP(clk), 
        .Q(n9628) );
  HS65_LS_DFPHQX4 clk_r_REG519_S1 ( .D(text_in_r[38]), .E(n9852), .CP(clk), 
        .Q(n9627) );
  HS65_LS_DFPHQX4 clk_r_REG520_S1 ( .D(text_in_r[37]), .E(n9852), .CP(clk), 
        .Q(n9626) );
  HS65_LS_DFPHQX4 clk_r_REG521_S1 ( .D(text_in_r[36]), .E(n9852), .CP(clk), 
        .Q(n9625) );
  HS65_LS_DFPHQX4 clk_r_REG522_S1 ( .D(text_in_r[35]), .E(n9852), .CP(clk), 
        .Q(n9624) );
  HS65_LS_DFPHQX4 clk_r_REG523_S1 ( .D(text_in_r[34]), .E(n9852), .CP(clk), 
        .Q(n9623) );
  HS65_LS_DFPHQX4 clk_r_REG524_S1 ( .D(text_in_r[33]), .E(n9852), .CP(clk), 
        .Q(n9622) );
  HS65_LS_DFPHQX4 clk_r_REG525_S1 ( .D(text_in_r[32]), .E(n9852), .CP(clk), 
        .Q(n9621) );
  HS65_LS_DFPHQX4 clk_r_REG526_S1 ( .D(text_in_r[31]), .E(n9852), .CP(clk), 
        .Q(n9620) );
  HS65_LS_DFPHQX4 clk_r_REG527_S1 ( .D(text_in_r[30]), .E(n9852), .CP(clk), 
        .Q(n9619) );
  HS65_LS_DFPHQX4 clk_r_REG528_S1 ( .D(text_in_r[29]), .E(n9851), .CP(clk), 
        .Q(n9618) );
  HS65_LS_DFPHQX4 clk_r_REG529_S1 ( .D(text_in_r[28]), .E(n9851), .CP(clk), 
        .Q(n9617) );
  HS65_LS_DFPHQX4 clk_r_REG530_S1 ( .D(text_in_r[27]), .E(n9851), .CP(clk), 
        .Q(n9616) );
  HS65_LS_DFPHQX4 clk_r_REG531_S1 ( .D(text_in_r[26]), .E(n9851), .CP(clk), 
        .Q(n9615) );
  HS65_LS_DFPHQX4 clk_r_REG532_S1 ( .D(text_in_r[25]), .E(n9851), .CP(clk), 
        .Q(n9614) );
  HS65_LS_DFPHQX4 clk_r_REG533_S1 ( .D(text_in_r[24]), .E(n9849), .CP(clk), 
        .Q(n9613) );
  HS65_LS_DFPHQX4 clk_r_REG534_S1 ( .D(text_in_r[23]), .E(n9851), .CP(clk), 
        .Q(n9612) );
  HS65_LS_DFPHQX4 clk_r_REG535_S1 ( .D(text_in_r[22]), .E(n9851), .CP(clk), 
        .Q(n9611) );
  HS65_LS_DFPHQX4 clk_r_REG536_S1 ( .D(text_in_r[21]), .E(n9851), .CP(clk), 
        .Q(n9610) );
  HS65_LS_DFPHQX4 clk_r_REG537_S1 ( .D(text_in_r[20]), .E(n9851), .CP(clk), 
        .Q(n9609) );
  HS65_LS_DFPHQX4 clk_r_REG538_S1 ( .D(text_in_r[19]), .E(n9851), .CP(clk), 
        .Q(n9608) );
  HS65_LS_DFPHQX4 clk_r_REG539_S1 ( .D(text_in_r[18]), .E(n9851), .CP(clk), 
        .Q(n9607) );
  HS65_LS_DFPHQX4 clk_r_REG540_S1 ( .D(text_in_r[17]), .E(n9851), .CP(clk), 
        .Q(n9606) );
  HS65_LS_DFPHQX4 clk_r_REG541_S1 ( .D(text_in_r[16]), .E(n9851), .CP(clk), 
        .Q(n9605) );
  HS65_LS_DFPHQX4 clk_r_REG542_S1 ( .D(text_in_r[15]), .E(n9851), .CP(clk), 
        .Q(n9604) );
  HS65_LS_DFPHQX4 clk_r_REG543_S1 ( .D(text_in_r[14]), .E(n9850), .CP(clk), 
        .Q(n9603) );
  HS65_LS_DFPHQX4 clk_r_REG544_S1 ( .D(text_in_r[13]), .E(n9850), .CP(clk), 
        .Q(n9602) );
  HS65_LS_DFPHQX4 clk_r_REG545_S1 ( .D(text_in_r[12]), .E(n9850), .CP(clk), 
        .Q(n9601) );
  HS65_LS_DFPHQX4 clk_r_REG546_S1 ( .D(text_in_r[11]), .E(n9850), .CP(clk), 
        .Q(n9600) );
  HS65_LS_DFPHQX4 clk_r_REG547_S1 ( .D(text_in_r[10]), .E(n9850), .CP(clk), 
        .Q(n9599) );
  HS65_LS_DFPHQX4 clk_r_REG548_S1 ( .D(text_in_r[9]), .E(n9850), .CP(clk), .Q(
        n9598) );
  HS65_LS_DFPHQX4 clk_r_REG549_S1 ( .D(text_in_r[8]), .E(n9850), .CP(clk), .Q(
        n9597) );
  HS65_LS_DFPHQX4 clk_r_REG550_S1 ( .D(text_in_r[7]), .E(n9850), .CP(clk), .Q(
        n9596) );
  HS65_LS_DFPHQX4 clk_r_REG551_S1 ( .D(text_in_r[6]), .E(n9850), .CP(clk), .Q(
        n9595) );
  HS65_LS_DFPHQX4 clk_r_REG552_S1 ( .D(text_in_r[5]), .E(n9850), .CP(clk), .Q(
        n9594) );
  HS65_LS_DFPHQX4 clk_r_REG553_S1 ( .D(text_in_r[4]), .E(n9850), .CP(clk), .Q(
        n9593) );
  HS65_LS_DFPHQX4 clk_r_REG554_S1 ( .D(text_in_r[3]), .E(n9850), .CP(clk), .Q(
        n9592) );
  HS65_LS_DFPHQX4 clk_r_REG555_S1 ( .D(text_in_r[2]), .E(n9850), .CP(clk), .Q(
        n9591) );
  HS65_LS_DFPHQX4 clk_r_REG556_S1 ( .D(text_in_r[1]), .E(n9850), .CP(clk), .Q(
        n9590) );
  HS65_LS_DFPHQX4 clk_r_REG557_S1 ( .D(text_in_r[0]), .E(n9849), .CP(clk), .Q(
        n9589) );
  HS65_LS_DFPQX4 clk_r_REG115_S6 ( .D(n2663), .CP(clk), .Q(n9456) );
  HS65_LS_DFPQX4 clk_r_REG167_S6 ( .D(n2747), .CP(clk), .Q(n9454) );
  HS65_LS_DFPQX4 clk_r_REG141_S23 ( .D(n5948), .CP(clk), .Q(n9424) );
  HS65_LS_DFPQX4 clk_r_REG135_S4 ( .D(n2751), .CP(clk), .Q(n9423) );
  HS65_LS_DFPQX4 clk_r_REG104_S9 ( .D(n7577), .CP(clk), .Q(n9422) );
  HS65_LS_DFPQX4 clk_r_REG145_S6 ( .D(n2625), .CP(clk), .Q(n9421) );
  HS65_LS_DFPQX4 clk_r_REG63_S16 ( .D(n4443), .CP(clk), .Q(n9420) );
  HS65_LS_DFPQX4 clk_r_REG41_S14 ( .D(n7605), .CP(clk), .Q(n9419) );
  HS65_LS_DFPQX4 clk_r_REG76_S14 ( .D(n2754), .CP(clk), .Q(n9418) );
  HS65_LS_DFPQX4 clk_r_REG101_S4 ( .D(n2742), .CP(clk), .Q(n9417) );
  HS65_LS_DFPQX4 clk_r_REG54_S16 ( .D(n2714), .CP(clk), .Q(n9416) );
  HS65_LS_DFPQX4 clk_r_REG129_S6 ( .D(n3546), .CP(clk), .Q(n9414) );
  HS65_LS_DFPQX4 clk_r_REG114_S14 ( .D(n7786), .CP(clk), .Q(n9413) );
  HS65_LS_DFPQX4 clk_r_REG50_S12 ( .D(n7608), .CP(clk), .Q(n9412) );
  HS65_LS_DFPQX4 clk_r_REG25_S5 ( .D(n7544), .CP(clk), .Q(n9411) );
  HS65_LS_DFPQX4 clk_r_REG56_S5 ( .D(sa02[7]), .CP(clk), .Q(n9403) );
  HS65_LS_DFPQX4 clk_r_REG170_S21 ( .D(sa00[7]), .CP(clk), .Q(n9402) );
  HS65_LS_DFPQX4 clk_r_REG158_S23 ( .D(sa31[3]), .CP(clk), .Q(n9401) );
  HS65_LS_DFPQX4 clk_r_REG178_S12 ( .D(sa20[5]), .CP(clk), .Q(n9399) );
  HS65_LS_DFPQX4 clk_r_REG200_S11 ( .D(sa01[2]), .CP(clk), .Q(n9396) );
  HS65_LS_DFPQX4 clk_r_REG156_S22 ( .D(sa01[0]), .CP(clk), .Q(n9392) );
  HS65_LS_DFPQX4 clk_r_REG47_S6 ( .D(sa12[7]), .CP(clk), .Q(n9390) );
  HS65_LS_DFPQX4 clk_r_REG212_S18 ( .D(sa11[6]), .CP(clk), .Q(n9389) );
  HS65_LS_DFPQX4 clk_r_REG187_S13 ( .D(sa10[6]), .CP(clk), .Q(n9388) );
  HS65_LS_DFPQX4 clk_r_REG57_S6 ( .D(sa32[5]), .CP(clk), .Q(n9387) );
  HS65_LS_DFPQX4 clk_r_REG189_S5 ( .D(sa11[7]), .CP(clk), .Q(n9385) );
  HS65_LS_DFPQX4 clk_r_REG190_S10 ( .D(sa20[0]), .CP(clk), .Q(n9384) );
  HS65_LS_DFPQX4 clk_r_REG133_S11 ( .D(sa10[7]), .CP(clk), .Q(n9383) );
  HS65_LS_DFPQX4 clk_r_REG148_S5 ( .D(sa31[7]), .CP(clk), .Q(n9382) );
  HS65_LS_DFPQX4 clk_r_REG161_S15 ( .D(sa30[7]), .CP(clk), .Q(n9381) );
  HS65_LS_DFPQX4 clk_r_REG168_S7 ( .D(sa11[0]), .CP(clk), .Q(n9380) );
  HS65_LS_DFPQX4 clk_r_REG86_S15 ( .D(sa22[0]), .CP(clk), .Q(n9379) );
  HS65_LS_DFPQX4 clk_r_REG163_S5 ( .D(sa21[0]), .CP(clk), .Q(n9378) );
  HS65_LS_DFPQX4 clk_r_REG30_S6 ( .D(sa32[2]), .CP(clk), .Q(n9377) );
  HS65_LS_DFPQX4 clk_r_REG73_S23 ( .D(sa31[2]), .CP(clk), .Q(n9376) );
  HS65_LS_DFPQX4 clk_r_REG81_S21 ( .D(sa30[6]), .CP(clk), .Q(n9374) );
  HS65_LS_DFPQX4 clk_r_REG107_S23 ( .D(sa31[6]), .CP(clk), .Q(n9373) );
  HS65_LS_DFPQX4 clk_r_REG98_S13 ( .D(sa30[0]), .CP(clk), .Q(n9372) );
  HS65_LS_DFPQX4 clk_r_REG16_S11 ( .D(sa31[0]), .CP(clk), .Q(n9371) );
  HS65_LS_DFPQX4 clk_r_REG108_S24 ( .D(sa02[0]), .CP(clk), .Q(n9370) );
  HS65_LS_DFPQX4 clk_r_REG37_S11 ( .D(sa30[2]), .CP(clk), .Q(n9369) );
  HS65_LS_DFPQX4 clk_r_REG10_S5 ( .D(sa32[6]), .CP(clk), .Q(n9368) );
  HS65_LS_DFPQX4 clk_r_REG93_S9 ( .D(sa30[5]), .CP(clk), .Q(n9367) );
  HS65_LS_DFPQX4 clk_r_REG109_S7 ( .D(sa32[4]), .CP(clk), .Q(n9366) );
  HS65_LS_DFPQX4 clk_r_REG82_S22 ( .D(sa21[6]), .CP(clk), .Q(n9365) );
  HS65_LS_DFPQX4 clk_r_REG18_S12 ( .D(sa22[5]), .CP(clk), .Q(n9364) );
  HS65_LS_DFPQX4 clk_r_REG159_S17 ( .D(sa22[4]), .CP(clk), .Q(n9362) );
  HS65_LS_DFPQX4 clk_r_REG125_S5 ( .D(sa32[3]), .CP(clk), .Q(n9361) );
  HS65_LS_DFPQX4 clk_r_REG49_S11 ( .D(sa31[1]), .CP(clk), .Q(n9360) );
  HS65_LS_DFPQX4 clk_r_REG59_S7 ( .D(sa21[2]), .CP(clk), .Q(n9358) );
  HS65_LS_DFPQX4 clk_r_REG123_S4 ( .D(sa02[4]), .CP(clk), .Q(n9356) );
  HS65_LS_DFPQX4 clk_r_REG99_S22 ( .D(sa21[4]), .CP(clk), .Q(n9355) );
  HS65_LS_DFPQX4 clk_r_REG102_S15 ( .D(sa11[3]), .CP(clk), .Q(n9354) );
  HS65_LS_DFPQX4 clk_r_REG48_S7 ( .D(sa01[3]), .CP(clk), .Q(n9353) );
  HS65_LS_DFPQX4 clk_r_REG149_S24 ( .D(sa22[3]), .CP(clk), .Q(n9352) );
  HS65_LS_DFPQX4 clk_r_REG62_S15 ( .D(sa22[1]), .CP(clk), .Q(n9351) );
  HS65_LS_DFPQX4 clk_r_REG22_S3 ( .D(sa21[1]), .CP(clk), .Q(n9350) );
  HS65_LS_DFPQX4 clk_r_REG95_S11 ( .D(sa11[1]), .CP(clk), .Q(n9349) );
  HS65_LS_DFPQX4 clk_r_REG143_S13 ( .D(sa31[4]), .CP(clk), .Q(n9348) );
  HS65_LS_DFPQX4 clk_r_REG138_S12 ( .D(sa20[4]), .CP(clk), .Q(n9347) );
  HS65_LS_DFPQX4 clk_r_REG77_S15 ( .D(sa11[4]), .CP(clk), .Q(n9346) );
  HS65_LS_DFPQX4 clk_r_REG21_S2 ( .D(sa12[4]), .CP(clk), .Q(n9345) );
  HS65_LS_DFPQX4 clk_r_REG27_S6 ( .D(sa02[1]), .CP(clk), .Q(n9344) );
  HS65_LS_DFPQX4 clk_r_REG13_S8 ( .D(sa20[3]), .CP(clk), .Q(n9342) );
  HS65_LS_DFPQX4 clk_r_REG120_S10 ( .D(sa21[3]), .CP(clk), .Q(n9341) );
  HS65_LS_DFPQX4 clk_r_REG75_S16 ( .D(sa10[4]), .CP(clk), .Q(n9340) );
  HS65_LS_DFPQX4 clk_r_REG45_S15 ( .D(sa02[3]), .CP(clk), .Q(n9336) );
  HS65_LS_DFPQX4 clk_r_REG140_S13 ( .D(sa12[5]), .CP(clk), .Q(n9335) );
  HS65_LS_DFPQX4 clk_r_REG31_S7 ( .D(sa03[1]), .CP(clk), .Q(n9334) );
  HS65_LS_DFPQX4 clk_r_REG97_S12 ( .D(sa00[1]), .CP(clk), .Q(n9333) );
  HS65_LS_DFPQX4 clk_r_REG15_S10 ( .D(sa01[1]), .CP(clk), .Q(n9332) );
  HS65_LS_DFPQX4 clk_r_REG172_S15 ( .D(sa10[0]), .CP(clk), .Q(n9330) );
  HS65_LS_DFPQX4 clk_r_REG113_S16 ( .D(sa20[6]), .CP(clk), .Q(n9329) );
  HS65_LS_DFPQX4 clk_r_REG71_S22 ( .D(sa01[4]), .CP(clk), .Q(n9328) );
  HS65_LS_DFPQX4 clk_r_REG87_S16 ( .D(sa10[3]), .CP(clk), .Q(n9327) );
  HS65_LS_DFPQX4 clk_r_REG136_S5 ( .D(sa11[2]), .CP(clk), .Q(n9325) );
  HS65_LS_DFPQX4 clk_r_REG150_S16 ( .D(sa10[2]), .CP(clk), .Q(n9324) );
  HS65_LS_DFPQX4 clk_r_REG103_S16 ( .D(sa20[2]), .CP(clk), .Q(n9322) );
  HS65_LS_DFPQX4 clk_r_REG69_S20 ( .D(sa00[3]), .CP(clk), .Q(n9321) );
  HS65_LS_DFPQX4 clk_r_REG35_S10 ( .D(sa00[4]), .CP(clk), .Q(n9320) );
  HS65_LS_DFPQX4 clk_r_REG183_S13 ( .D(sa12[0]), .CP(clk), .Q(n9318) );
  HS65_LS_DFPQX4 clk_r_REG126_S7 ( .D(sa03[0]), .CP(clk), .Q(n9316) );
  HS65_LS_DFPQX4 clk_r_REG127_S8 ( .D(sa13[7]), .CP(clk), .Q(n9314) );
  HS65_LS_DFPQX4 clk_r_REG121_S8 ( .D(sa13[6]), .CP(clk), .Q(n9313) );
  HS65_LS_DFPQX4 clk_r_REG118_S10 ( .D(sa00[0]), .CP(clk), .Q(n9312) );
  HS65_LS_DFPQX4 clk_r_REG165_S17 ( .D(sa03[4]), .CP(clk), .Q(n9310) );
  HS65_LS_DFPQX4 clk_r_REG111_S8 ( .D(sa23[6]), .CP(clk), .Q(n9308) );
  HS65_LS_DFPQX4 clk_r_REG33_S9 ( .D(sa33[1]), .CP(clk), .Q(n9307) );
  HS65_LS_DFPQX4 clk_r_REG12_S7 ( .D(sa33[4]), .CP(clk), .Q(n9306) );
  HS65_LS_DFPQX4 clk_r_REG58_S6 ( .D(sa23[7]), .CP(clk), .Q(n9305) );
  HS65_LS_DFPQX4 clk_r_REG67_S19 ( .D(sa33[7]), .CP(clk), .Q(n9302) );
  HS65_LS_DFPQX4 clk_r_REG52_S14 ( .D(sa23[0]), .CP(clk), .Q(n9301) );
  HS65_LS_DFPQX4 clk_r_REG32_S8 ( .D(sa03[7]), .CP(clk), .Q(n9299) );
  HS65_LS_DFPQX4 clk_r_REG44_S14 ( .D(sa13[3]), .CP(clk), .Q(n9247) );
  HS65_LS_DFPQX4 clk_r_REG19_S13 ( .D(sa20[7]), .CP(clk), .Q(n9246) );
  HS65_LS_DFPQX4 clk_r_REG7_S3 ( .D(sa13[4]), .CP(clk), .Q(n9245) );
  HS65_LS_DFPQX4 clk_r_REG119_S13 ( .D(sa30[4]), .CP(clk), .Q(n9244) );
  HS65_LS_DFPQX4 clk_r_REG28_S5 ( .D(sa02[2]), .CP(clk), .Q(n9243) );
  HS65_LS_DFPQX4 clk_r_REG70_S21 ( .D(sa30[1]), .CP(clk), .Q(n9242) );
  HS65_LS_DFPQX4 clk_r_REG23_S4 ( .D(sa13[1]), .CP(clk), .Q(n9241) );
  HS65_LS_DFPQX4 clk_r_REG64_S17 ( .D(sa12[3]), .CP(clk), .Q(n9240) );
  HS65_LS_DFPQX4 clk_r_REG14_S9 ( .D(sa12[1]), .CP(clk), .Q(n9239) );
  HS65_LS_DFPQX4 clk_r_REG51_S13 ( .D(sa10[1]), .CP(clk), .Q(n9238) );
  HS65_LS_DFPQX4 clk_r_REG155_S11 ( .D(sa30[3]), .CP(clk), .Q(n9237) );
  HS65_LS_DFPQX4 clk_r_REG91_S8 ( .D(sa00[6]), .CP(clk), .Q(n9236) );
  HS65_LS_DFPQX4 clk_r_REG38_S12 ( .D(sa01[6]), .CP(clk), .Q(n9235) );
  HS65_LS_DFPQX4 clk_r_REG324_S6 ( .D(w3[18]), .CP(clk), .Q(n9174) );
  HS65_LS_DFPQX4 clk_r_REG312_S7 ( .D(w3[26]), .CP(clk), .Q(n9169) );
  HS65_LS_DFPQNX4 clk_r_REG371_S8 ( .D(\u0/N46 ), .CP(clk), .QN(n954) );
  HS65_LS_DFPQNX4 clk_r_REG342_S8 ( .D(\u0/N45 ), .CP(clk), .QN(n953) );
  HS65_LS_BFX2 U9543 ( .A(n9859), .Z(n9861) );
  HS65_LS_BFX2 U9544 ( .A(n9866), .Z(n9859) );
  HS65_LS_IVX4 U9545 ( .A(n9859), .Z(n9853) );
  HS65_LS_IVX2 U9546 ( .A(ld), .Z(n9866) );
  HS65_LS_BFX4 U9547 ( .A(n9866), .Z(n9860) );
  HS65_LS_IVX4 U9548 ( .A(n9860), .Z(n9857) );
  HS65_LS_IVX4 U9549 ( .A(n9860), .Z(n9858) );
  HS65_LS_BFX2 U9550 ( .A(n9860), .Z(n9865) );
  HS65_LS_IVX2 U9551 ( .A(n9860), .Z(n9846) );
  HS65_LS_IVX4 U9552 ( .A(n9860), .Z(n9847) );
  HS65_LS_IVX4 U9647 ( .A(n9860), .Z(n9848) );
  HS65_LS_IVX4 U9648 ( .A(n9861), .Z(n9849) );
  HS65_LS_IVX4 U9649 ( .A(n9860), .Z(n9850) );
  HS65_LS_IVX4 U9650 ( .A(n9860), .Z(n9851) );
  HS65_LS_IVX4 U9651 ( .A(n9860), .Z(n9852) );
  HS65_LS_IVX4 U9652 ( .A(n9860), .Z(n9854) );
  HS65_LS_IVX2 U13189 ( .A(n9860), .Z(n9855) );
  HS65_LS_IVX2 U13200 ( .A(n9860), .Z(n9856) );
  HS65_LS_BFX2 U13201 ( .A(n9861), .Z(n9862) );
  HS65_LS_BFX4 U13206 ( .A(n9859), .Z(n9863) );
  HS65_LS_BFX4 U16895 ( .A(n9865), .Z(n9864) );
  HS65_LS_DFPQX4 clk_r_REG293_S7 ( .D(n7576), .CP(clk), .Q(n9477) );
  HS65_LS_DFPQX4 clk_r_REG399_S9 ( .D(n2624), .CP(clk), .Q(n9476) );
  HS65_LS_DFPQX4 clk_r_REG318_S6 ( .D(n4442), .CP(clk), .Q(n9475) );
  HS65_LS_DFPQX4 clk_r_REG391_S10 ( .D(n7607), .CP(clk), .Q(n9435) );
  HS65_LS_DFPQX4 clk_r_REG276_S6 ( .D(n7604), .CP(clk), .Q(n9474) );
  HS65_LS_DFPQX4 clk_r_REG297_S8 ( .D(n5947), .CP(clk), .Q(n9570) );
  HS65_LS_DFPQX4 clk_r_REG404_S5 ( .D(n7785), .CP(clk), .Q(n9436) );
  HS65_LS_DFPQX4 clk_r_REG380_S8 ( .D(n7543), .CP(clk), .Q(n9434) );
  HS65_LS_DFPQX4 clk_r_REG321_S6 ( .D(n2753), .CP(clk), .Q(n9461) );
  HS65_LS_DFPQX4 clk_r_REG362_S10 ( .D(n2741), .CP(clk), .Q(n9460) );
  HS65_LS_DFPQX4 clk_r_REG401_S6 ( .D(n2750), .CP(clk), .Q(n9569) );
  HS65_LS_DFPQX4 clk_r_REG313_S8 ( .D(n2670), .CP(clk), .Q(n9458) );
  HS65_LS_DFPQX4 clk_r_REG325_S7 ( .D(n2713), .CP(clk), .Q(n9459) );
  HS65_LS_DFPQX4 clk_r_REG349_S10 ( .D(n2746), .CP(clk), .Q(n9455) );
  HS65_LS_DFPQX4 clk_r_REG345_S9 ( .D(n3545), .CP(clk), .Q(n9437) );
  HS65_LS_DFPQX4 clk_r_REG341_S4 ( .D(n2662), .CP(clk), .Q(n9457) );
  HS65_LS_DFPQX4 clk_r_REG418_S2 ( .D(n9148), .CP(clk), .Q(n9575) );
  HS65_LS_DFPQX4 clk_r_REG420_S2 ( .D(n9147), .CP(clk), .Q(n9578) );
  HS65_LS_DFPQX4 clk_r_REG419_S2 ( .D(n9142), .CP(clk), .Q(n9582) );
  HS65_LS_DFPQX4 clk_r_REG426_S2 ( .D(n9140), .CP(clk), .Q(n9587) );
  HS65_LS_DFPQX4 clk_r_REG423_S2 ( .D(n9144), .CP(clk), .Q(n9581) );
  HS65_LS_DFPQX4 clk_r_REG424_S2 ( .D(n9138), .CP(clk), .Q(n9584) );
  HS65_LS_DFPQX4 clk_r_REG427_S2 ( .D(n9141), .CP(clk), .Q(n9585) );
  HS65_LS_DFPQX4 clk_r_REG425_S2 ( .D(n9139), .CP(clk), .Q(n9586) );
  HS65_LS_DFPQX4 clk_r_REG422_S2 ( .D(n9143), .CP(clk), .Q(n9580) );
  HS65_LS_DFPQX4 clk_r_REG421_S2 ( .D(n9145), .CP(clk), .Q(n9576) );
  HS65_LS_DFPQX4 clk_r_REG429_S1 ( .D(\u0/r0/rcnt [1]), .CP(clk), .Q(n9579) );
  HS65_LS_DFPQX4 clk_r_REG415_S2 ( .D(\u0/rcon [24]), .CP(clk), .Q(n9163) );
  HS65_LS_DFPQX4 clk_r_REG428_S1 ( .D(\u0/r0/rcnt [0]), .CP(clk), .Q(n9577) );
  HS65_LS_DFPQX4 clk_r_REG3_S1 ( .D(dcnt[2]), .CP(clk), .Q(n9407) );
  HS65_LS_DFPQX4 clk_r_REG417_S1 ( .D(n9858), .CP(clk), .Q(n9588) );
  HS65_LS_DFPQX4 clk_r_REG407_S1 ( .D(\u0/r0/rcnt [3]), .CP(clk), .Q(n9571) );
  HS65_LS_DFPQX4 clk_r_REG412_S2 ( .D(\u0/rcon [27]), .CP(clk), .Q(n9162) );
  HS65_LS_DFPQX4 clk_r_REG1_S1 ( .D(dcnt[3]), .CP(clk), .Q(n9164) );
  HS65_LS_DFPQX4 clk_r_REG4_S1 ( .D(dcnt[0]), .CP(clk), .Q(n9408) );
  HS65_LS_DFPQX4 clk_r_REG416_S1 ( .D(\u0/r0/rcnt [2]), .CP(clk), .Q(n9572) );
  HS65_LS_DFPQX4 clk_r_REG0_S1 ( .D(dcnt[1]), .CP(clk), .Q(n9161) );
  HS65_LS_DFPQX4 clk_r_REG413_S2 ( .D(\u0/rcon [26]), .CP(clk), .Q(n9404) );
  HS65_LS_DFPQX4 clk_r_REG228_S14 ( .D(n629), .CP(clk), .Q(n9583) );
  HS65_LS_DFPQX4 clk_r_REG414_S2 ( .D(\u0/rcon [25]), .CP(clk), .Q(n9406) );
  HS65_LS_DFPQX4 clk_r_REG408_S2 ( .D(\u0/rcon [31]), .CP(clk), .Q(n9410) );
  HS65_LS_DFPQX4 clk_r_REG410_S2 ( .D(\u0/rcon [30]), .CP(clk), .Q(n9425) );
  HS65_LS_DFPQX4 clk_r_REG411_S2 ( .D(\u0/rcon [28]), .CP(clk), .Q(n9405) );
  HS65_LS_DFPQX4 clk_r_REG409_S2 ( .D(\u0/rcon [29]), .CP(clk), .Q(n9165) );
  HS65_LS_DFPQX4 clk_r_REG269_S4 ( .D(w0[5]), .CP(clk), .Q(n9226) );
  HS65_LS_DFPQX4 clk_r_REG302_S9 ( .D(w0[13]), .CP(clk), .Q(n9215) );
  HS65_LS_DFPQX4 clk_r_REG284_S4 ( .D(w0[7]), .CP(clk), .Q(n9263) );
  HS65_LS_DFPQX4 clk_r_REG335_S6 ( .D(w0[21]), .CP(clk), .Q(n9199) );
  HS65_LS_DFPQX4 clk_r_REG273_S5 ( .D(w0[15]), .CP(clk), .Q(n9266) );
  HS65_LS_DFPQX4 clk_r_REG317_S5 ( .D(w0[9]), .CP(clk), .Q(n9264) );
  HS65_LS_DFPQX4 clk_r_REG374_S9 ( .D(w0[8]), .CP(clk), .Q(n9258) );
  HS65_LS_DFPQX4 clk_r_REG306_S10 ( .D(w0[23]), .CP(clk), .Q(n9261) );
  HS65_LS_DFPQX4 clk_r_REG278_S6 ( .D(w0[17]), .CP(clk), .Q(n9267) );
  HS65_LS_DFPQX4 clk_r_REG365_S6 ( .D(w0[16]), .CP(clk), .Q(n9259) );
  HS65_LS_DFPQX4 clk_r_REG314_S8 ( .D(w0[6]), .CP(clk), .Q(n9268) );
  HS65_LS_DFPQX4 clk_r_REG359_S9 ( .D(w0[12]), .CP(clk), .Q(n9214) );
  HS65_LS_DFPQX4 clk_r_REG363_S6 ( .D(w0[20]), .CP(clk), .Q(n9211) );
  HS65_LS_DFPQX4 clk_r_REG346_S9 ( .D(w0[11]), .CP(clk), .Q(n9269) );
  HS65_LS_DFPQX4 clk_r_REG290_S6 ( .D(w0[22]), .CP(clk), .Q(n9271) );
  HS65_LS_DFPQX4 clk_r_REG332_S9 ( .D(w0[14]), .CP(clk), .Q(n9273) );
  HS65_LS_DFPQX4 clk_r_REG329_S8 ( .D(w0[0]), .CP(clk), .Q(n9257) );
  HS65_LS_DFPQX4 clk_r_REG299_S8 ( .D(w0[1]), .CP(clk), .Q(n9272) );
  HS65_LS_DFPQX4 clk_r_REG281_S7 ( .D(w0[29]), .CP(clk), .Q(n9194) );
  HS65_LS_DFPQX4 clk_r_REG350_S6 ( .D(w0[19]), .CP(clk), .Q(n9270) );
  HS65_LS_DFPQX4 clk_r_REG270_S4 ( .D(w1[5]), .CP(clk), .Q(n9212) );
  HS65_LS_DFPQX4 clk_r_REG295_S7 ( .D(w0[31]), .CP(clk), .Q(n9248) );
  HS65_LS_DFPQX4 clk_r_REG303_S9 ( .D(w1[13]), .CP(clk), .Q(n9209) );
  HS65_LS_DFPQX4 clk_r_REG265_S3 ( .D(w0[25]), .CP(clk), .Q(n9262) );
  HS65_LS_DFPQX4 clk_r_REG353_S3 ( .D(w0[24]), .CP(clk), .Q(n9260) );
  HS65_LS_DFPQX4 clk_r_REG336_S6 ( .D(w1[21]), .CP(clk), .Q(n9202) );
  HS65_LS_DFPQX4 clk_r_REG326_S7 ( .D(w0[28]), .CP(clk), .Q(n9193) );
  HS65_LS_DFPQX4 clk_r_REG285_S4 ( .D(w1[7]), .CP(clk), .Q(n9229) );
  HS65_LS_DFPQX4 clk_r_REG368_S7 ( .D(w0[30]), .CP(clk), .Q(n9331) );
  HS65_LS_DFPQX4 clk_r_REG330_S8 ( .D(w1[0]), .CP(clk), .Q(n9228) );
  HS65_LS_DFPQX4 clk_r_REG338_S3 ( .D(w0[27]), .CP(clk), .Q(n9265) );
  HS65_LS_DFPQX4 clk_r_REG300_S8 ( .D(w1[1]), .CP(clk), .Q(n9223) );
  HS65_LS_DFPQX4 clk_r_REG356_S4 ( .D(w0[2]), .CP(clk), .Q(n9225) );
  HS65_LS_DFPQX4 clk_r_REG319_S5 ( .D(w1[9]), .CP(clk), .Q(n9221) );
  HS65_LS_DFPQX4 clk_r_REG274_S5 ( .D(w1[15]), .CP(clk), .Q(n9217) );
  HS65_LS_DFPQX4 clk_r_REG360_S9 ( .D(w1[12]), .CP(clk), .Q(n9208) );
  HS65_LS_DFPQX4 clk_r_REG307_S10 ( .D(w1[23]), .CP(clk), .Q(n9231) );
  HS65_LS_DFPQX4 clk_r_REG375_S9 ( .D(w1[8]), .CP(clk), .Q(n9232) );
  HS65_LS_DFPQX4 clk_r_REG372_S8 ( .D(w1[4]), .CP(clk), .Q(n9207) );
  HS65_LS_DFPQX4 clk_r_REG279_S6 ( .D(w1[17]), .CP(clk), .Q(n9219) );
  HS65_LS_DFPQX4 clk_r_REG287_S5 ( .D(w0[10]), .CP(clk), .Q(n9196) );
  HS65_LS_DFPQX4 clk_r_REG315_S8 ( .D(w1[6]), .CP(clk), .Q(n9227) );
  HS65_LS_DFPQX4 clk_r_REG366_S6 ( .D(w1[16]), .CP(clk), .Q(n9230) );
  HS65_LS_DFPQX4 clk_r_REG364_S6 ( .D(w1[20]), .CP(clk), .Q(n9206) );
  HS65_LS_DFPQX4 clk_r_REG322_S6 ( .D(w0[18]), .CP(clk), .Q(n9195) );
  HS65_LS_DFPQX4 clk_r_REG201_S16 ( .D(n2673), .CP(clk), .Q(n9574) );
  HS65_LS_DFPQX4 clk_r_REG282_S7 ( .D(w1[29]), .CP(clk), .Q(n9200) );
  HS65_LS_DFPQX4 clk_r_REG333_S9 ( .D(w1[14]), .CP(clk), .Q(n9224) );
  HS65_LS_DFPQX4 clk_r_REG343_S8 ( .D(w1[3]), .CP(clk), .Q(n9222) );
  HS65_LS_DFPQX4 clk_r_REG271_S4 ( .D(w2[5]), .CP(clk), .Q(n9287) );
  HS65_LS_DFPQX4 clk_r_REG347_S9 ( .D(w1[11]), .CP(clk), .Q(n9216) );
  HS65_LS_DFPQX4 clk_r_REG291_S6 ( .D(w1[22]), .CP(clk), .Q(n9233) );
  HS65_LS_DFPQX4 clk_r_REG304_S9 ( .D(w2[13]), .CP(clk), .Q(n9286) );
  HS65_LS_DFPQX4 clk_r_REG351_S6 ( .D(w1[19]), .CP(clk), .Q(n9218) );
  HS65_LS_DFPQX4 clk_r_REG296_S7 ( .D(w1[31]), .CP(clk), .Q(n9205) );
  HS65_LS_DFPQX4 clk_r_REG389_S6 ( .D(w2[21]), .CP(clk), .Q(n9249) );
  HS65_LS_DFPQX4 clk_r_REG403_S4 ( .D(w2[7]), .CP(clk), .Q(n9294) );
  HS65_LS_DFPQX4 clk_r_REG266_S3 ( .D(w1[25]), .CP(clk), .Q(n9204) );
  HS65_LS_DFPQX4 clk_r_REG354_S3 ( .D(w1[24]), .CP(clk), .Q(n9234) );
  HS65_LS_DFPQX4 clk_r_REG327_S7 ( .D(w1[28]), .CP(clk), .Q(n9197) );
  HS65_LS_DFPQX4 clk_r_REG392_S8 ( .D(w2[0]), .CP(clk), .Q(n9282) );
  HS65_LS_DFPQX4 clk_r_REG398_S8 ( .D(w2[1]), .CP(clk), .Q(n9285) );
  HS65_LS_DFPQX4 clk_r_REG275_S5 ( .D(w2[15]), .CP(clk), .Q(n9254) );
  HS65_LS_DFPQX4 clk_r_REG395_S5 ( .D(w2[9]), .CP(clk), .Q(n9293) );
  HS65_LS_DFPQX4 clk_r_REG310_S7 ( .D(w0[26]), .CP(clk), .Q(n9192) );
  HS65_LS_DFPQX4 clk_r_REG377_S9 ( .D(w2[8]), .CP(clk), .Q(n9297) );
  HS65_LS_DFPQX4 clk_r_REG308_S1 ( .D(w2[23]), .CP(clk), .Q(n9280) );
  HS65_LS_DFPQX4 clk_r_REG357_S4 ( .D(w1[2]), .CP(clk), .Q(n9213) );
  HS65_LS_DFPQX4 clk_r_REG396_S8 ( .D(w2[6]), .CP(clk), .Q(n9291) );
  HS65_LS_DFPQX4 clk_r_REG369_S7 ( .D(w1[30]), .CP(clk), .Q(n9203) );
  HS65_LS_DFPQX4 clk_r_REG378_S1 ( .D(w2[4]), .CP(clk), .Q(n9289) );
  HS65_LS_DFPQX4 clk_r_REG382_S9 ( .D(w2[12]), .CP(clk), .Q(n9288) );
  HS65_LS_DFPQX4 clk_r_REG381_S6 ( .D(w2[16]), .CP(clk), .Q(n9256) );
  HS65_LS_DFPQX4 clk_r_REG339_S3 ( .D(w1[27]), .CP(clk), .Q(n9220) );
  HS65_LS_DFPQX4 clk_r_REG406_S1 ( .D(w2[17]), .CP(clk), .Q(n9253) );
  HS65_LS_DFPQX4 clk_r_REG405_S1 ( .D(w2[29]), .CP(clk), .Q(n9275) );
  HS65_LS_DFPQX4 clk_r_REG390_S9 ( .D(w2[14]), .CP(clk), .Q(n9284) );
  HS65_LS_DFPQX4 clk_r_REG5_S1 ( .D(w2[20]), .CP(clk), .Q(n9251) );
  HS65_LS_DFPQX4 clk_r_REG387_S8 ( .D(w2[3]), .CP(clk), .Q(n9296) );
  HS65_LS_DFPQX4 clk_r_REG386_S9 ( .D(w2[11]), .CP(clk), .Q(n9290) );
  HS65_LS_DFPQX4 clk_r_REG292_S6 ( .D(w2[22]), .CP(clk), .Q(n9250) );
  HS65_LS_DFPQX4 clk_r_REG288_S5 ( .D(w1[10]), .CP(clk), .Q(n9210) );
  HS65_LS_DFPQX4 clk_r_REG272_S4 ( .D(w3[5]), .CP(clk), .Q(n9393) );
  HS65_LS_DFPQX4 clk_r_REG323_S6 ( .D(w1[18]), .CP(clk), .Q(n9201) );
  HS65_LS_DFPQX4 clk_r_REG305_S9 ( .D(w3[13]), .CP(clk), .Q(n9339) );
  HS65_LS_DFPQX4 clk_r_REG385_S6 ( .D(w2[19]), .CP(clk), .Q(n9252) );
  HS65_LS_DFPQX4 clk_r_REG90_S9 ( .D(sa33[5]), .CP(clk), .Q(n9311) );
  HS65_LS_DFPQX4 clk_r_REG400_S7 ( .D(w2[31]), .CP(clk), .Q(n9283) );
  HS65_LS_DFPQX4 clk_r_REG393_S7 ( .D(w2[28]), .CP(clk), .Q(n9276) );
  HS65_LS_DFPQX4 clk_r_REG267_S3 ( .D(w2[25]), .CP(clk), .Q(n9279) );
  HS65_LS_DFPQX4 clk_r_REG384_S3 ( .D(w2[24]), .CP(clk), .Q(n9281) );
  HS65_LS_DFPQX4 clk_r_REG337_S6 ( .D(w3[21]), .CP(clk), .Q(n9172) );
  HS65_LS_DFPQX4 clk_r_REG286_S4 ( .D(w3[7]), .CP(clk), .Q(n9171) );
  HS65_LS_DFPQX4 clk_r_REG331_S8 ( .D(w3[0]), .CP(clk), .Q(n9191) );
  HS65_LS_DFPQX4 clk_r_REG152_S17 ( .D(sa03[5]), .CP(clk), .Q(n9315) );
  HS65_LS_DFPQX4 clk_r_REG131_S13 ( .D(sa00[5]), .CP(clk), .Q(n9400) );
  HS65_LS_DFPQX4 clk_r_REG301_S8 ( .D(w3[1]), .CP(clk), .Q(n9178) );
  HS65_LS_DFPQX4 clk_r_REG320_S5 ( .D(w3[9]), .CP(clk), .Q(n9176) );
  HS65_LS_DFPQX4 clk_r_REG277_S5 ( .D(w3[15]), .CP(clk), .Q(n9338) );
  HS65_LS_DFPQX4 clk_r_REG376_S9 ( .D(w3[8]), .CP(clk), .Q(n9189) );
  HS65_LS_DFPQX4 clk_r_REG309_S10 ( .D(w3[23]), .CP(clk), .Q(n9386) );
  HS65_LS_DFPQX4 clk_r_REG311_S7 ( .D(w1[26]), .CP(clk), .Q(n9198) );
  HS65_LS_DFPQX4 clk_r_REG361_S9 ( .D(w3[12]), .CP(clk), .Q(n9185) );
  HS65_LS_DFPQX4 clk_r_REG383_S4 ( .D(w2[2]), .CP(clk), .Q(n9292) );
  HS65_LS_DFPQX4 clk_r_REG379_S7 ( .D(w2[30]), .CP(clk), .Q(n9274) );
  HS65_LS_DFPQX4 clk_r_REG316_S8 ( .D(w3[6]), .CP(clk), .Q(n9188) );
  HS65_LS_DFPQX4 clk_r_REG373_S8 ( .D(w3[4]), .CP(clk), .Q(n9186) );
  HS65_LS_DFPQX4 clk_r_REG106_S22 ( .D(sa01[5]), .CP(clk), .Q(n9395) );
  HS65_LS_DFPQX4 clk_r_REG147_S17 ( .D(sa23[5]), .CP(clk), .Q(n9398) );
  HS65_LS_DFPQX4 clk_r_REG83_S16 ( .D(sa13[5]), .CP(clk), .Q(n9309) );
  HS65_LS_DFPQX4 clk_r_REG89_S17 ( .D(sa03[6]), .CP(clk), .Q(n9298) );
  HS65_LS_DFPQX4 clk_r_REG283_S7 ( .D(w3[29]), .CP(clk), .Q(n9181) );
  HS65_LS_DFPQX4 clk_r_REG280_S6 ( .D(w3[17]), .CP(clk), .Q(n9167) );
  HS65_LS_DFPQX4 clk_r_REG367_S6 ( .D(w3[16]), .CP(clk), .Q(n9173) );
  HS65_LS_DFPQX4 clk_r_REG6_S2 ( .D(w3[20]), .CP(clk), .Q(n9175) );
  HS65_LS_DFPQX4 clk_r_REG388_S3 ( .D(w2[27]), .CP(clk), .Q(n9278) );
  HS65_LS_DFPQX4 clk_r_REG334_S9 ( .D(w3[14]), .CP(clk), .Q(n9182) );
  HS65_LS_DFPQX4 clk_r_REG344_S8 ( .D(w3[3]), .CP(clk), .Q(n9180) );
  HS65_LS_DFPQX4 clk_r_REG348_S9 ( .D(w3[11]), .CP(clk), .Q(n9177) );
  HS65_LS_DFPQX4 clk_r_REG402_S5 ( .D(w2[10]), .CP(clk), .Q(n9295) );
  HS65_LS_DFPQX4 clk_r_REG294_S6 ( .D(w3[22]), .CP(clk), .Q(n9394) );
  HS65_LS_DFPQX4 clk_r_REG40_S13 ( .D(sa31[5]), .CP(clk), .Q(n9375) );
  HS65_LS_DFPQX4 clk_r_REG394_S1 ( .D(w2[18]), .CP(clk), .Q(n9255) );
  HS65_LS_DFPQX4 clk_r_REG74_S15 ( .D(sa22[2]), .CP(clk), .Q(n9363) );
  HS65_LS_DFPQX4 clk_r_REG53_S15 ( .D(sa21[7]), .CP(clk), .Q(n9343) );
  HS65_LS_DFPQX4 clk_r_REG8_S4 ( .D(sa02[5]), .CP(clk), .Q(n9357) );
  HS65_LS_DFPQX4 clk_r_REG298_S7 ( .D(w3[31]), .CP(clk), .Q(n9183) );
  HS65_LS_DFPQX4 clk_r_REG352_S6 ( .D(w3[19]), .CP(clk), .Q(n9168) );
  HS65_LS_DFPQX4 clk_r_REG328_S7 ( .D(w3[28]), .CP(clk), .Q(n9179) );
  HS65_LS_DFPQX4 clk_r_REG268_S3 ( .D(w3[25]), .CP(clk), .Q(n9337) );
  HS65_LS_DFPQX4 clk_r_REG355_S3 ( .D(w3[24]), .CP(clk), .Q(n9187) );
  HS65_LS_DFPQX4 clk_r_REG42_S13 ( .D(sa10[5]), .CP(clk), .Q(n9323) );
  HS65_LS_DFPQX4 clk_r_REG79_S21 ( .D(sa00[2]), .CP(clk), .Q(n9397) );
  HS65_LS_DFPQX4 clk_r_REG179_S13 ( .D(sa12[2]), .CP(clk), .Q(n9303) );
  HS65_LS_DFPQX4 clk_r_REG11_S6 ( .D(n2672), .CP(clk), .Q(n9415) );
  HS65_LS_DFPQX4 clk_r_REG397_S1 ( .D(w2[26]), .CP(clk), .Q(n9277) );
  HS65_LS_DFPQX4 clk_r_REG175_S8 ( .D(sa33[6]), .CP(clk), .Q(n9319) );
  HS65_LS_DFPQX4 clk_r_REG370_S7 ( .D(w3[30]), .CP(clk), .Q(n9170) );
  HS65_LS_DFPQX4 clk_r_REG358_S4 ( .D(w3[2]), .CP(clk), .Q(n9190) );
  HS65_LS_DFPQX4 clk_r_REG153_S6 ( .D(sa33[0]), .CP(clk), .Q(n9300) );
  HS65_LS_DFPQX4 clk_r_REG340_S3 ( .D(w3[27]), .CP(clk), .Q(n9166) );
  HS65_LS_DFPQX4 clk_r_REG116_S7 ( .D(sa33[2]), .CP(clk), .Q(n9304) );
  HS65_LS_DFPQX4 clk_r_REG185_S6 ( .D(sa32[0]), .CP(clk), .Q(n9391) );
  HS65_LS_DFPQX4 clk_r_REG289_S5 ( .D(w3[10]), .CP(clk), .Q(n9184) );
  HS65_LS_DFPQX4 clk_r_REG66_S18 ( .D(sa21[5]), .CP(clk), .Q(n9359) );
  HS65_LS_DFPQX4 clk_r_REG112_S7 ( .D(sa11[5]), .CP(clk), .Q(n9326) );
  HS65_LS_DFPQX4 clk_r_REG60_S14 ( .D(sa13[0]), .CP(clk), .Q(n9317) );
  HS65_LSS_DFPQX18 clk_r_REG2_S2 ( .D(n9717), .CP(clk), .Q(done) );
  HS65_LSS_DFPQX18 clk_r_REG206_S10 ( .D(n9749), .CP(clk), .Q(text_out[96]) );
  HS65_LSS_DFPQX18 clk_r_REG263_S6 ( .D(n9843), .CP(clk), .Q(text_out[2]) );
  HS65_LSS_DFPQX18 clk_r_REG254_S5 ( .D(n9788), .CP(clk), .Q(text_out[57]) );
  HS65_LSS_DFPQX18 clk_r_REG117_S8 ( .D(n9748), .CP(clk), .Q(text_out[97]) );
  HS65_LSS_DFPQX18 clk_r_REG216_S9 ( .D(n9799), .CP(clk), .Q(text_out[46]) );
  HS65_LSS_DFPQX18 clk_r_REG84_S15 ( .D(n9791), .CP(clk), .Q(text_out[54]) );
  HS65_LSS_DFPQX18 clk_r_REG198_S3 ( .D(n9759), .CP(clk), .Q(text_out[86]) );
  HS65_LSS_DFPQX18 clk_r_REG221_S8 ( .D(n9743), .CP(clk), .Q(text_out[102]) );
  HS65_LSS_DFPQX18 clk_r_REG249_S14 ( .D(n9807), .CP(clk), .Q(text_out[38]) );
  HS65_LSS_DFPQX18 clk_r_REG245_S11 ( .D(n9756), .CP(clk), .Q(text_out[89]) );
  HS65_LSS_DFPQX18 clk_r_REG151_S3 ( .D(n9825), .CP(clk), .Q(text_out[20]) );
  HS65_LSS_DFPQX18 clk_r_REG193_S22 ( .D(n9781), .CP(clk), .Q(text_out[64]) );
  HS65_LSS_DFPQX18 clk_r_REG188_S7 ( .D(n9773), .CP(clk), .Q(text_out[72]) );
  HS65_LSS_DFPQX18 clk_r_REG207_S7 ( .D(n9819), .CP(clk), .Q(text_out[26]) );
  HS65_LSS_DFPQX18 clk_r_REG34_S10 ( .D(n9745), .CP(clk), .Q(text_out[100]) );
  HS65_LSS_DFPQX18 clk_r_REG256_S3 ( .D(n9764), .CP(clk), .Q(text_out[81]) );
  HS65_LSS_DFPQX18 clk_r_REG237_S7 ( .D(n9772), .CP(clk), .Q(text_out[73]) );
  HS65_LSS_DFPQX18 clk_r_REG239_S6 ( .D(n9784), .CP(clk), .Q(text_out[61]) );
  HS65_LSS_DFPQX18 clk_r_REG252_S8 ( .D(n9815), .CP(clk), .Q(text_out[30]) );
  HS65_LSS_DFPQX18 clk_r_REG68_S20 ( .D(n9746), .CP(clk), .Q(text_out[99]) );
  HS65_LSS_DFPQX18 clk_r_REG166_S9 ( .D(n9818), .CP(clk), .Q(text_out[27]) );
  HS65_LSS_DFPQX18 clk_r_REG243_S13 ( .D(n9740), .CP(clk), .Q(text_out[105])
         );
  HS65_LSS_DFPQX18 clk_r_REG213_S7 ( .D(n9785), .CP(clk), .Q(text_out[60]) );
  HS65_LSS_DFPQX18 clk_r_REG218_S15 ( .D(n9770), .CP(clk), .Q(text_out[75]) );
  HS65_LSS_DFPQX18 clk_r_REG259_S10 ( .D(n9765), .CP(clk), .Q(text_out[80]) );
  HS65_LSS_DFPQX18 clk_r_REG258_S11 ( .D(n9757), .CP(clk), .Q(text_out[88]) );
  HS65_LSS_DFPQX18 clk_r_REG235_S16 ( .D(n9741), .CP(clk), .Q(text_out[104])
         );
  HS65_LSS_DFPQX18 clk_r_REG9_S5 ( .D(n9783), .CP(clk), .Q(text_out[62]) );
  HS65_LSS_DFPQX18 clk_r_REG241_S15 ( .D(n9767), .CP(clk), .Q(text_out[78]) );
  HS65_LSS_DFPQX18 clk_r_REG210_S16 ( .D(n9727), .CP(clk), .Q(text_out[118])
         );
  HS65_LSS_DFPQX18 clk_r_REG238_S6 ( .D(n9838), .CP(clk), .Q(text_out[7]) );
  HS65_LSS_DFPQX18 clk_r_REG215_S23 ( .D(n9751), .CP(clk), .Q(text_out[94]) );
  HS65_LSS_DFPQX18 clk_r_REG226_S15 ( .D(n9769), .CP(clk), .Q(text_out[76]) );
  HS65_LSS_DFPQX18 clk_r_REG194_S18 ( .D(n9821), .CP(clk), .Q(text_out[24]) );
  HS65_LSS_DFPQX18 clk_r_REG55_S15 ( .D(n9790), .CP(clk), .Q(text_out[55]) );
  HS65_LSS_DFPQX18 clk_r_REG17_S12 ( .D(n9809), .CP(clk), .Q(text_out[36]) );
  HS65_LSS_DFPQX18 clk_r_REG224_S16 ( .D(n9832), .CP(clk), .Q(text_out[13]) );
  HS65_LSS_DFPQX18 clk_r_REG88_S17 ( .D(n9824), .CP(clk), .Q(text_out[21]) );
  HS65_LSS_DFPQX18 clk_r_REG164_S8 ( .D(n9833), .CP(clk), .Q(text_out[12]) );
  HS65_LSS_DFPQX18 clk_r_REG169_S12 ( .D(n9726), .CP(clk), .Q(text_out[119])
         );
  HS65_LSS_DFPQX18 clk_r_REG137_S12 ( .D(n9729), .CP(clk), .Q(text_out[116])
         );
  HS65_LSS_DFPQX18 clk_r_REG227_S14 ( .D(n9828), .CP(clk), .Q(text_out[17]) );
  HS65_LSS_DFPQX18 clk_r_REG196_S24 ( .D(n9811), .CP(clk), .Q(text_out[34]) );
  HS65_LSS_DFPQX18 clk_r_REG177_S12 ( .D(n9728), .CP(clk), .Q(text_out[117])
         );
  HS65_LSS_DFPQX18 clk_r_REG205_S13 ( .D(n9721), .CP(clk), .Q(text_out[124])
         );
  HS65_LSS_DFPQX18 clk_r_REG139_S13 ( .D(n9800), .CP(clk), .Q(text_out[45]) );
  HS65_LSS_DFPQX18 clk_r_REG176_S12 ( .D(n9730), .CP(clk), .Q(text_out[115])
         );
  HS65_LSS_DFPQX18 clk_r_REG171_S9 ( .D(n9722), .CP(clk), .Q(text_out[123]) );
  HS65_LSS_DFPQX18 clk_r_REG92_S9 ( .D(n9720), .CP(clk), .Q(text_out[125]) );
  HS65_LSS_DFPQX18 clk_r_REG174_S17 ( .D(n9823), .CP(clk), .Q(text_out[22]) );
  HS65_LSS_DFPQX18 clk_r_REG225_S22 ( .D(n9776), .CP(clk), .Q(text_out[69]) );
  HS65_LSS_DFPQX18 clk_r_REG242_S14 ( .D(n9829), .CP(clk), .Q(text_out[16]) );
  HS65_LSS_DFPQX18 clk_r_REG217_S16 ( .D(n9731), .CP(clk), .Q(text_out[114])
         );
  HS65_LSS_DFPQX18 clk_r_REG162_S12 ( .D(n9774), .CP(clk), .Q(text_out[71]) );
  HS65_LSS_DFPQX18 clk_r_REG36_S11 ( .D(n9723), .CP(clk), .Q(text_out[122]) );
  HS65_LSS_DFPQX18 clk_r_REG132_S11 ( .D(n9718), .CP(clk), .Q(text_out[127])
         );
  HS65_LSS_DFPQX18 clk_r_REG186_S7 ( .D(n9840), .CP(clk), .Q(text_out[5]) );
  HS65_LSS_DFPQX18 clk_r_REG144_S14 ( .D(n9806), .CP(clk), .Q(text_out[39]) );
  HS65_LSS_DFPQX18 clk_r_REG204_S10 ( .D(n9779), .CP(clk), .Q(text_out[66]) );
  HS65_LSS_DFPQX18 clk_r_REG146_S7 ( .D(n9841), .CP(clk), .Q(text_out[4]) );
  HS65_LSS_DFPQX18 clk_r_REG20_S14 ( .D(n9801), .CP(clk), .Q(text_out[44]) );
  HS65_LSS_DFPQX18 clk_r_REG173_S17 ( .D(n9826), .CP(clk), .Q(text_out[19]) );
  HS65_LSS_DFPQX18 clk_r_REG24_S5 ( .D(n9792), .CP(clk), .Q(text_out[53]) );
  HS65_LSS_DFPQX18 clk_r_REG46_S6 ( .D(n9782), .CP(clk), .Q(text_out[63]) );
  HS65_LSS_DFPQX18 clk_r_REG236_S8 ( .D(n9837), .CP(clk), .Q(text_out[8]) );
  HS65_LSS_DFPQX18 clk_r_REG255_S4 ( .D(n9836), .CP(clk), .Q(text_out[9]) );
  HS65_LSS_DFPQX18 clk_r_REG248_S13 ( .D(n9736), .CP(clk), .Q(text_out[109])
         );
  HS65_LSS_DFPQX18 clk_r_REG180_S10 ( .D(n9758), .CP(clk), .Q(text_out[87]) );
  HS65_LSS_DFPQX18 clk_r_REG195_S16 ( .D(n9739), .CP(clk), .Q(text_out[106])
         );
  HS65_LSS_DFPQX18 clk_r_REG105_S7 ( .D(n9761), .CP(clk), .Q(text_out[84]) );
  HS65_LSS_DFPQX18 clk_r_REG182_S13 ( .D(n9803), .CP(clk), .Q(text_out[42]) );
  HS65_LSS_DFPQX18 clk_r_REG203_S8 ( .D(n9831), .CP(clk), .Q(text_out[14]) );
  HS65_LSS_DFPQX18 clk_r_REG43_S14 ( .D(n9822), .CP(clk), .Q(text_out[23]) );
  HS65_LSS_DFPQX18 clk_r_REG191_S24 ( .D(n9810), .CP(clk), .Q(text_out[35]) );
  HS65_LSS_DFPQX18 clk_r_REG100_S4 ( .D(n9834), .CP(clk), .Q(text_out[11]) );
  HS65_LSS_DFPQX18 clk_r_REG65_S18 ( .D(n9760), .CP(clk), .Q(text_out[85]) );
  HS65_LSS_DFPQX18 clk_r_REG39_S13 ( .D(n9752), .CP(clk), .Q(text_out[93]) );
  HS65_LSS_DFPQX18 clk_r_REG262_S7 ( .D(n9817), .CP(clk), .Q(text_out[28]) );
  HS65_LSS_DFPQX18 clk_r_REG233_S19 ( .D(n9830), .CP(clk), .Q(text_out[15]) );
  HS65_LSS_DFPQX18 clk_r_REG29_S6 ( .D(n9787), .CP(clk), .Q(text_out[58]) );
  HS65_LSS_DFPQX18 clk_r_REG181_S18 ( .D(n9762), .CP(clk), .Q(text_out[83]) );
  HS65_LSS_DFPQX18 clk_r_REG211_S7 ( .D(n9768), .CP(clk), .Q(text_out[77]) );
  HS65_LSS_DFPQX18 clk_r_REG247_S15 ( .D(n9795), .CP(clk), .Q(text_out[50]) );
  HS65_LSS_DFPQX18 clk_r_REG72_S23 ( .D(n9755), .CP(clk), .Q(text_out[90]) );
  HS65_LSS_DFPQX18 clk_r_REG192_S13 ( .D(n9750), .CP(clk), .Q(text_out[95]) );
  HS65_LSS_DFPQX18 clk_r_REG157_S23 ( .D(n9754), .CP(clk), .Q(text_out[91]) );
  HS65_LSS_DFPQX18 clk_r_REG230_S24 ( .D(n9812), .CP(clk), .Q(text_out[33]) );
  HS65_LSS_DFPQX18 clk_r_REG142_S13 ( .D(n9753), .CP(clk), .Q(text_out[92]) );
  HS65_LSS_DFPQX18 clk_r_REG222_S9 ( .D(n9816), .CP(clk), .Q(text_out[29]) );
  HS65_LSS_DFPQX18 clk_r_REG122_S4 ( .D(n9794), .CP(clk), .Q(text_out[51]) );
  HS65_LSS_DFPQX18 clk_r_REG80_S21 ( .D(n9719), .CP(clk), .Q(text_out[126]) );
  HS65_LSS_DFPQX18 clk_r_REG199_S5 ( .D(n9771), .CP(clk), .Q(text_out[74]) );
  HS65_LSS_DFPQX18 clk_r_REG154_S10 ( .D(n9742), .CP(clk), .Q(text_out[103])
         );
  HS65_LSS_DFPQX18 clk_r_REG244_S12 ( .D(n9808), .CP(clk), .Q(text_out[37]) );
  HS65_LSS_DFPQX18 clk_r_REG246_S7 ( .D(n9763), .CP(clk), .Q(text_out[82]) );
  HS65_LSS_DFPQX18 clk_r_REG160_S15 ( .D(n9734), .CP(clk), .Q(text_out[111])
         );
  HS65_LSS_DFPQX18 clk_r_REG209_S14 ( .D(n9798), .CP(clk), .Q(text_out[47]) );
  HS65_LSS_DFPQX18 clk_r_REG130_S10 ( .D(n9744), .CP(clk), .Q(text_out[101])
         );
  HS65_LSS_DFPQX18 clk_r_REG96_S12 ( .D(n9733), .CP(clk), .Q(text_out[112]) );
  HS65_LSS_DFPQX18 clk_r_REG234_S17 ( .D(n9802), .CP(clk), .Q(text_out[43]) );
  HS65_LSS_DFPQX18 clk_r_REG26_S6 ( .D(n9789), .CP(clk), .Q(text_out[56]) );
  HS65_LSS_DFPQX18 clk_r_REG202_S7 ( .D(n9845), .CP(clk), .Q(text_out[0]) );
  HS65_LSS_DFPQX18 clk_r_REG220_S13 ( .D(n9725), .CP(clk), .Q(text_out[120])
         );
  HS65_LSS_DFPQX18 clk_r_REG219_S22 ( .D(n9778), .CP(clk), .Q(text_out[67]) );
  HS65_LSS_DFPQX18 clk_r_REG253_S7 ( .D(n9844), .CP(clk), .Q(text_out[1]) );
  HS65_LSS_DFPQX18 clk_r_REG231_S22 ( .D(n9777), .CP(clk), .Q(text_out[68]) );
  HS65_LSS_DFPQX18 clk_r_REG240_S16 ( .D(n9835), .CP(clk), .Q(text_out[10]) );
  HS65_LSS_DFPQX18 clk_r_REG264_S2 ( .D(n9793), .CP(clk), .Q(text_out[52]) );
  HS65_LSS_DFPQX18 clk_r_REG251_S9 ( .D(n9820), .CP(clk), .Q(text_out[25]) );
  HS65_LSS_DFPQX18 clk_r_REG261_S8 ( .D(n9747), .CP(clk), .Q(text_out[98]) );
  HS65_LSS_DFPQX18 clk_r_REG197_S5 ( .D(n9766), .CP(clk), .Q(text_out[79]) );
  HS65_LSS_DFPQX18 clk_r_REG110_S7 ( .D(n9839), .CP(clk), .Q(text_out[6]) );
  HS65_LSS_DFPQX18 clk_r_REG134_S17 ( .D(n9827), .CP(clk), .Q(text_out[18]) );
  HS65_LSS_DFPQX18 clk_r_REG78_S16 ( .D(n9732), .CP(clk), .Q(text_out[113]) );
  HS65_LSS_DFPQX18 clk_r_REG85_S15 ( .D(n9797), .CP(clk), .Q(text_out[48]) );
  HS65_LSS_DFPQX18 clk_r_REG208_S6 ( .D(n9842), .CP(clk), .Q(text_out[3]) );
  HS65_LSS_DFPQX18 clk_r_REG229_S16 ( .D(n9737), .CP(clk), .Q(text_out[108])
         );
  HS65_LSS_DFPQX18 clk_r_REG61_S15 ( .D(n9796), .CP(clk), .Q(text_out[49]) );
  HS65_LSS_DFPQX18 clk_r_REG124_S5 ( .D(n9786), .CP(clk), .Q(text_out[59]) );
  HS65_LSS_DFPQX18 clk_r_REG257_S13 ( .D(n9735), .CP(clk), .Q(text_out[110])
         );
  HS65_LSS_DFPQX18 clk_r_REG232_S21 ( .D(n9724), .CP(clk), .Q(text_out[121])
         );
  HS65_LSS_DFPQX18 clk_r_REG128_S8 ( .D(n9814), .CP(clk), .Q(text_out[31]) );
  HS65_LSS_DFPQX18 clk_r_REG214_S24 ( .D(n9813), .CP(clk), .Q(text_out[32]) );
  HS65_LSS_DFPQX18 clk_r_REG223_S16 ( .D(n9738), .CP(clk), .Q(text_out[107])
         );
  HS65_LSS_DFPQX18 clk_r_REG260_S9 ( .D(n9804), .CP(clk), .Q(text_out[41]) );
  HS65_LSS_DFPQX18 clk_r_REG184_S13 ( .D(n9805), .CP(clk), .Q(text_out[40]) );
  HS65_LSS_DFPQX18 clk_r_REG94_S10 ( .D(n9780), .CP(clk), .Q(text_out[65]) );
  HS65_LSS_DFPQX18 clk_r_REG250_S12 ( .D(n9775), .CP(clk), .Q(text_out[70]) );
endmodule

